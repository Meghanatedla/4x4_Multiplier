*** 4 BIT MULTIPLIER

.INCLUDE ../TSMC_180nm.txt

.INCLUDE AND.sub
.INCLUDE HA.sub
.INCLUDE FA.sub

*PARAMETERS
.PARAM X=0.09u

.PARAM Width_p=10*X
.PARAM Length_p=2*X

.PARAM Width_n=5*X
.PARAM Length_n=2*X

.PARAM supply=1
.PARAM tr=10p

.global gnd vdd

.temp 25

*NET-LIST

* Inputs: A3 A2 A1 A0   B3 B2 B1 B0
* Outputs: C S6 S5 S4 S3 S2 S1 S0
* 16 AND gates
* 4 Half adders
* 8 Full adders
* Inputs nodes to HA  is given as HA_ax HA_bx (x = 1, 2, 3, 4)
* Inputs nodes to FA  is given as FA_ax FA_bx FA_cx (x = 1, 2, 3, 4, 5, 6, 7, 8)

xAnd1   A0 B0 vdd gnd  S0   AND
xAnd2   A0 B1 vdd gnd HA_a1 AND
xAnd3   A1 B0 vdd gnd HA_b1 AND
xAnd4   A0 B2 vdd gnd FA_a1 AND
xAnd5   A2 B0 vdd gnd HA_a2 AND
xAnd6   A1 B1 vdd gnd HA_b2 AND
xAnd7   A1 B2 vdd gnd FA_a3 AND
xAnd8   A0 B3 vdd gnd FA_b2 AND
xAnd9   A3 B0 vdd gnd HA_a4 AND
xAnd10  A2 B1 vdd gnd HA_b4 AND
xAnd11  A2 B2 vdd gnd FA_a7 AND
xAnd12  A3 B1 vdd gnd FA_b7 AND
xAnd13  A1 B3 vdd gnd FA_b4 AND
xAnd14  A2 B3 vdd gnd FA_a8 AND
xAnd15  A3 B2 vdd gnd FA_b8 AND
xAnd16  A3 B3 vdd gnd FA_b6 AND

xHA1 HA_a1 HA_b1 vdd gnd  S1   FA_c1 HA
xHA2 HA_a2 HA_b2 vdd gnd FA_b1 FA_c3 HA
xHA3 HA_a3 HA_b3 vdd gnd  S4   FA_c5 HA
xHA4 HA_a4 HA_b4 vdd gnd FA_b3 FA_c7 HA

xFA1 FA_a1 FA_b1 FA_c1 vdd gnd  S2   FA_c2 FA
xFA2 FA_a2 FA_b2 FA_c2 vdd gnd  S3   HA_a3 FA
xFA3 FA_a3 FA_b3 FA_c3 vdd gnd FA_a2 FA_c4 FA
xFA4 FA_a4 FA_b4 FA_c4 vdd gnd HA_b3 FA_a5 FA
xFA5 FA_a5 FA_b5 FA_c5 vdd gnd  S5   FA_c6 FA
xFA6 FA_a6 FA_b6 FA_c6 vdd gnd  S6     C   FA
xFA7 FA_a7 FA_b7 FA_c7 vdd gnd FA_a4 FA_c8 FA
xFA8 FA_a8 FA_b8 FA_c8 vdd gnd FA_b5 FA_a6 FA

*SOURCE
VDD vdd gnd 'supply'

*Capacitive LOAD
CL1 S0 gnd 0.01f
CL2 S1 gnd 0.01f
CL3 S2 gnd 0.01f
CL4 S3 gnd 0.01f
CL5 S4 gnd 0.01f
CL6 S5 gnd 0.01f
CL7 S6 gnd 0.01f
CL8 C  gnd 0.01f

*INPUT WAVEFORM
VA0 A0 gnd PWL(0 0 {0+500m} 0 {0+500m+tr} 1 {0+1000m} 1 {0+1000m+tr} 0 {0+1500m} 0 {0+1500m+tr} 1 {0+2000m} 1 {0+2000m+tr} 0 {0+2500m} 0 {0+2500m+tr} 1 {0+3000m} 1 {0+3000m+tr} 0 {0+3500m} 0 {0+3500m+tr} 1 {0+4000m} 1 {0+4000m+tr} 0 {0+4500m} 0 {0+4500m+tr} 1 {0+5000m} 1 {0+5000m+tr} 0 {0+5500m} 0 {0+5500m+tr} 1 {0+6000m} 1 {0+6000m+tr} 0 {0+6500m} 0 {0+6500m+tr} 1 {0+7000m} 1 {0+7000m+tr} 0 {0+7500m} 0 {0+7500m+tr} 1 {0+8000m} 1 {0+8000m+tr} 0 {0+8500m} 0 {0+8500m+tr} 1 {0+9000m} 1 {0+9000m+tr} 1 {0+9500m} 1 {0+9500m+tr} 0)
VA1 A1 gnd PWL(0 0 {0+500m} 0 {0+500m+tr} 0 {0+1000m} 0 {0+1000m+tr} 1 {0+1500m} 1 {0+1500m+tr} 1 {0+2000m} 1 {0+2000m+tr} 0 {0+2500m} 0 {0+2500m+tr} 0 {0+3000m} 0 {0+3000m+tr} 1 {0+3500m} 1 {0+3500m+tr} 1 {0+4000m} 1 {0+4000m+tr} 0 {0+4500m} 0 {0+4500m+tr} 0 {0+5000m} 0 {0+5000m+tr} 1 {0+5500m} 1 {0+5500m+tr} 1 {0+6000m} 1 {0+6000m+tr} 0 {0+6500m} 0 {0+6500m+tr} 0 {0+7000m} 0 {0+7000m+tr} 0 {0+7500m} 0 {0+7500m+tr} 1 {0+8000m} 1 {0+8000m+tr} 1 {0+8500m} 1 {0+8500m+tr} 0 {0+9000m} 0 {0+9000m+tr} 0 {0+9500m} 0 {0+9500m+tr} 1)
VA2 A2 gnd PWL(0 0 {0+500m} 0 {0+500m+tr} 0 {0+1000m} 0 {0+1000m+tr} 0 {0+1500m} 0 {0+1500m+tr} 0 {0+2000m} 0 {0+2000m+tr} 1 {0+2500m} 1 {0+2500m+tr} 1 {0+3000m} 1 {0+3000m+tr} 1 {0+3500m} 1 {0+3500m+tr} 1 {0+4000m} 1 {0+4000m+tr} 0 {0+4500m} 0 {0+4500m+tr} 0 {0+5000m} 0 {0+5000m+tr} 1 {0+5500m} 1 {0+5500m+tr} 1 {0+6000m} 1 {0+6000m+tr} 0 {0+6500m} 0 {0+6500m+tr} 1 {0+7000m} 1 {0+7000m+tr} 1 {0+7500m} 1 {0+7500m+tr} 1 {0+8000m} 1 {0+8000m+tr} 0 {0+8500m} 0 {0+8500m+tr} 1 {0+9000m} 1 {0+9000m+tr} 1 {0+9500m} 1 {0+9500m+tr} 0)
VA3 A3 gnd PWL(0 0 {0+500m} 0 {0+500m+tr} 0 {0+1000m} 0 {0+1000m+tr} 0 {0+1500m} 0 {0+1500m+tr} 0 {0+2000m} 0 {0+2000m+tr} 1 {0+2500m} 1 {0+2500m+tr} 1 {0+3000m} 1 {0+3000m+tr} 1 {0+3500m} 1 {0+3500m+tr} 1 {0+4000m} 1 {0+4000m+tr} 0 {0+4500m} 0 {0+4500m+tr} 0 {0+5000m} 0 {0+5000m+tr} 1 {0+5500m} 1 {0+5500m+tr} 1 {0+6000m} 1 {0+6000m+tr} 1 {0+6500m} 1 {0+6500m+tr} 1 {0+7000m} 1 {0+7000m+tr} 1 {0+7500m} 1 {0+7500m+tr} 1 {0+8000m} 1 {0+8000m+tr} 1 {0+8500m} 1 {0+8500m+tr} 1 {0+9000m} 1 {0+9000m+tr} 1 {0+9500m} 1 {0+9500m+tr} 1)

VB0 B0 gnd PWL(0 0 {0+500m} 0 {0+500m+tr} 1 {0+1000m} 1 {0+1000m+tr} 0 {0+1500m} 0 {0+1500m+tr} 1 {0+2000m} 1 {0+2000m+tr} 0 {0+2500m} 0 {0+2500m+tr} 1 {0+3000m} 1 {0+3000m+tr} 0 {0+3500m} 0 {0+3500m+tr} 1 {0+4000m} 1 {0+4000m+tr} 1 {0+4500m} 1 {0+4500m+tr} 0 {0+5000m} 0 {0+5000m+tr} 1 {0+5500m} 1 {0+5500m+tr} 0 {0+6000m} 0 {0+6000m+tr} 0 {0+6500m} 0 {0+6500m+tr} 1 {0+7000m} 1 {0+7000m+tr} 1 {0+7500m} 1 {0+7500m+tr} 0 {0+8000m} 0 {0+8000m+tr} 0 {0+8500m} 0 {0+8500m+tr} 1 {0+9000m} 1 {0+9000m+tr} 0 {0+9500m} 0 {0+9500m+tr} 1)
VB1 B1 gnd PWL(0 0 {0+500m} 0 {0+500m+tr} 0 {0+1000m} 0 {0+1000m+tr} 1 {0+1500m} 1 {0+1500m+tr} 1 {0+2000m} 1 {0+2000m+tr} 0 {0+2500m} 0 {0+2500m+tr} 0 {0+3000m} 0 {0+3000m+tr} 1 {0+3500m} 1 {0+3500m+tr} 1 {0+4000m} 1 {0+4000m+tr} 1 {0+4500m} 1 {0+4500m+tr} 1 {0+5000m} 1 {0+5000m+tr} 0 {0+5500m} 0 {0+5500m+tr} 0 {0+6000m} 0 {0+6000m+tr} 0 {0+6500m} 0 {0+6500m+tr} 0 {0+7000m} 0 {0+7000m+tr} 0 {0+7500m} 0 {0+7500m+tr} 1 {0+8000m} 1 {0+8000m+tr} 1 {0+8500m} 1 {0+8500m+tr} 0 {0+9000m} 0 {0+9000m+tr} 1 {0+9500m} 1 {0+9500m+tr} 0)
VB2 B2 gnd PWL(0 0 {0+500m} 0 {0+500m+tr} 0 {0+1000m} 0 {0+1000m+tr} 0 {0+1500m} 0 {0+1500m+tr} 0 {0+2000m} 0 {0+2000m+tr} 1 {0+2500m} 1 {0+2500m+tr} 1 {0+3000m} 1 {0+3000m+tr} 1 {0+3500m} 1 {0+3500m+tr} 1 {0+4000m} 1 {0+4000m+tr} 1 {0+4500m} 1 {0+4500m+tr} 1 {0+5000m} 1 {0+5000m+tr} 0 {0+5500m} 0 {0+5500m+tr} 0 {0+6000m} 0 {0+6000m+tr} 1 {0+6500m} 1 {0+6500m+tr} 1 {0+7000m} 1 {0+7000m+tr} 1 {0+7500m} 1 {0+7500m+tr} 1 {0+8000m} 1 {0+8000m+tr} 0 {0+8500m} 0 {0+8500m+tr} 0 {0+9000m} 0 {0+9000m+tr} 0 {0+9500m} 0 {0+9500m+tr} 0)
VB3 B3 gnd PWL(0 0 {0+500m} 0 {0+500m+tr} 0 {0+1000m} 0 {0+1000m+tr} 0 {0+1500m} 0 {0+1500m+tr} 0 {0+2000m} 0 {0+2000m+tr} 1 {0+2500m} 1 {0+2500m+tr} 1 {0+3000m} 1 {0+3000m+tr} 1 {0+3500m} 1 {0+3500m+tr} 1 {0+4000m} 1 {0+4000m+tr} 1 {0+4500m} 1 {0+4500m+tr} 1 {0+5000m} 1 {0+5000m+tr} 0 {0+5500m} 0 {0+5500m+tr} 0 {0+6000m} 0 {0+6000m+tr} 1 {0+6500m} 1 {0+6500m+tr} 0 {0+7000m} 0 {0+7000m+tr} 1 {0+7500m} 1 {0+7500m+tr} 1 {0+8000m} 1 {0+8000m+tr} 0 {0+8500m} 0 {0+8500m+tr} 1 {0+9000m} 1 {0+9000m+tr} 1 {0+9500m} 1 {0+9500m+tr} 1)


*ANALYSIS
.TRAN 0.1m {10000m}

.CONTROL
set hcopypscolor = 1 
set color0=white 
set color1=black 

run

*******************************************
* A0
meas tran delay_LH_A0_S0
+ TRIG v(A0) val = 0.5 rise = 1
+ TARG v(S0) val = 0.5 rise = 1
meas tran delay_HL_A0_S0
+ TRIG v(A0) val = 0.5 fall = 1
+ TARG v(S0) val = 0.5 fall = 1
let delay_A0_S0 = (delay_LH_A0_S0+delay_HL_A0_S0)/2

meas tran delay_LH_A0_S1
+ TRIG v(A0) val = 0.5 rise = 5
+ TARG v(S1) val = 0.5 rise = 3
meas tran delay_HL_A0_S1
+ TRIG v(A0) val = 0.5 rise = 6
+ TARG v(S1) val = 0.5 fall = 3
let delay_A0_S1 = (delay_LH_A0_S1+delay_HL_A0_S1)/2

meas tran delay_LH_A0_S2
+ TRIG v(A0) val = 0.5 fall = 1
+ TARG v(S2) val = 0.5 rise = 1
meas tran delay_HL_A0_S2
+ TRIG v(A0) val = 0.5 rise = 2
+ TARG v(S2) val = 0.5 fall = 1
let delay_A0_S2 = (delay_LH_A0_S2+delay_HL_A0_S2)/2

meas tran delay_LH_A0_S3
+ TRIG v(A0) val = 0.5 fall = 7
+ TARG v(S3) val = 0.5 rise = 6
meas tran delay_HL_A0_S3
+ TRIG v(A0) val = 0.5 rise = 6
+ TARG v(S3) val = 0.5 fall = 5
let delay_A0_S3 = (delay_LH_A0_S3+delay_HL_A0_S3)/2

meas tran delay_LH_A0_S4
+ TRIG v(A0) val = 0.5 fall = 2
+ TARG v(S4) val = 0.5 rise = 1
meas tran delay_HL_A0_S4
+ TRIG v(A0) val = 0.5 rise = 3
+ TARG v(S4) val = 0.5 fall = 1
let delay_A0_S4 = (delay_LH_A0_S4+delay_HL_A0_S4)/2

meas tran delay_LH_A0_S5
+ TRIG v(A0) val = 0.5 fall = 6
+ TARG v(S5) val = 0.5 rise = 3
meas tran delay_HL_A0_S5
+ TRIG v(A0) val = 0.5 rise = 7
+ TARG v(S5) val = 0.5 fall = 3
let delay_A0_S5 = (delay_LH_A0_S5+delay_HL_A0_S5)/2

meas tran delay_LH_A0_S6
+ TRIG v(A0) val = 0.5 fall = 3
+ TARG v(S6) val = 0.5 rise = 2
meas tran delay_HL_A0_S6
+ TRIG v(A0) val = 0.5 rise = 7
+ TARG v(S6) val = 0.5 fall = 3
let delay_A0_S6 = (delay_LH_A0_S6+delay_HL_A0_S6)/2

meas tran delay_LH_A0_C
+ TRIG v(A0) val = 0.5 fall = 2
+ TARG v(C) val = 0.5 rise = 1
meas tran delay_HL_A0_C
+ TRIG v(A0) val = 0.5 fall = 4
+ TARG v(C) val = 0.5 fall = 1 
let delay_A0_C = (delay_LH_A0_C+delay_HL_A0_C)/2 

echo "A0">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo "Delay_LH_A0_S0 = $&delay_LH_A0_S0">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_HL_A0_S0 = $&delay_HL_A0_S0">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_A0_S0 = $&delay_A0_S0" >> "4_bit_Multiplier_Pre_Layout_pd.txt"
echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo "Delay_LH_A0_S1 = $&delay_LH_A0_S1">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_HL_A0_S1 = $&delay_HL_A0_S1">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_A0_S1 = $&delay_A0_S1" >> "4_bit_Multiplier_Pre_Layout_pd.txt"
echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo "Delay_LH_A0_S2 = $&delay_LH_A0_S2">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_HL_A0_S2 = $&delay_HL_A0_S2">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_A0_S2 = $&delay_A0_S2" >> "4_bit_Multiplier_Pre_Layout_pd.txt"
echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo "Delay_LH_A0_S3 = $&delay_LH_A0_S3">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_HL_A0_S3 = $&delay_HL_A0_S3">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_A0_S3 = $&delay_A0_S3" >> "4_bit_Multiplier_Pre_Layout_pd.txt"
echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo "Delay_LH_A0_S4 = $&delay_LH_A0_S4">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_HL_A0_S4 = $&delay_HL_A0_S4">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_A0_S4 = $&delay_A0_S4" >> "4_bit_Multiplier_Pre_Layout_pd.txt"
echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo "Delay_LH_A0_S5 = $&delay_LH_A0_S5">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_HL_A0_S5 = $&delay_HL_A0_S5">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_A0_S5 = $&delay_A0_S5" >> "4_bit_Multiplier_Pre_Layout_pd.txt"
echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo "Delay_LH_A0_S6 = $&delay_LH_A0_S6">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_HL_A0_S6 = $&delay_HL_A0_S6">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_A0_S6 = $&delay_A0_S6" >> "4_bit_Multiplier_Pre_Layout_pd.txt"
echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo "Delay_LH_A0_C = $&delay_LH_A0_C">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_HL_A0_C = $&delay_HL_A0_C">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_A0_C = $&delay_A0_C" >> "4_bit_Multiplier_Pre_Layout_pd.txt"
echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

****************************************************

* A1
meas tran delay_LH_A1_S0
+ TRIG v(A1) val = 0.5 fall = 4
+ TARG v(S0) val = 0.5 rise = 6
meas tran delay_HL_A1_S0
+ TRIG v(A1) val = 0.5 rise = 1
+ TARG v(S0) val = 0.5 fall = 1
let delay_A1_S0 = (delay_LH_A1_S0+delay_HL_A1_S0)/2

meas tran delay_LH_A1_S2
+ TRIG v(A1) val = 0.5 rise = 1
+ TARG v(S2) val = 0.5 rise = 1
meas tran delay_HL_A1_S2
+ TRIG v(A1) val = 0.5 rise = 3
+ TARG v(S2) val = 0.5 fall = 4
let delay_A1_S2 = (delay_LH_A1_S2+delay_HL_A1_S2)/2

meas tran delay_LH_A1_S3
+ TRIG v(A1) val = 0.5 fall = 4
+ TARG v(S3) val = 0.5 rise = 7
meas tran delay_HL_A1_S3
+ TRIG v(A1) val = 0.5 rise = 2
+ TARG v(S3) val = 0.5 fall = 2
let delay_A1_S3 = (delay_LH_A1_S3+delay_HL_A1_S3)/2

meas tran delay_LH_A1_S4
+ TRIG v(A1) val = 0.5 fall = 1
+ TARG v(S4) val = 0.5 rise = 1
meas tran delay_HL_A1_S4
+ TRIG v(A1) val = 0.5 rise = 4
+ TARG v(S4) val = 0.5 fall = 4
let delay_A1_S4 = (delay_LH_A1_S4+delay_HL_A1_S4)/2

meas tran delay_LH_A1_S5 
+ TRIG v(A1) val = 0.5 fall = 3
+ TARG v(S5) val = 0.5 rise = 3
meas tran delay_HL_A1_S5
+ TRIG v(A1) val = 0.5 rise = 2
+ TARG v(S5) val = 0.5 fall = 1
let delay_A1_S5 = (delay_LH_A1_S5+delay_HL_A1_S5)/2

meas tran delay_LH_A1_S6
+ TRIG v(A1) val = 0.5 fall = 1
+ TARG v(S6) val = 0.5 rise = 1
meas tran delay_HL_A1_S6
+ TRIG v(A1) val = 0.5 fall = 2
+ TARG v(S6) val = 0.5 fall = 2
let delay_A1_S6 = (delay_LH_A1_S6+delay_HL_A1_S6)/2

meas tran delay_LH_A1_C
+ TRIG v(A1) val = 0.5 fall = 1
+ TARG v(C) val = 0.5 rise = 1
meas tran delay_HL_A1_C
+ TRIG v(A1) val = 0.5 rise = 5
+ TARG v(C) val = 0.5 fall = 3 
let delay_A1_C = (delay_LH_A1_C+delay_HL_A1_C)/2 

echo "A1">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo "Delay_LH_A1_S0 = $&delay_LH_A1_S0">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_HL_A1_S0 = $&delay_HL_A1_S0">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_A1_S0 = $&delay_A1_S0" >> "4_bit_Multiplier_Pre_Layout_pd.txt"
echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo "Delay_LH_A1_S2 = $&delay_LH_A1_S2">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_HL_A1_S2 = $&delay_HL_A1_S2">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_A1_S2 = $&delay_A1_S2" >> "4_bit_Multiplier_Pre_Layout_pd.txt"
echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo "Delay_LH_A1_S3 = $&delay_LH_A1_S3">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_HL_A1_S3 = $&delay_HL_A1_S3">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_A1_S3 = $&delay_A1_S3" >> "4_bit_Multiplier_Pre_Layout_pd.txt"
echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo "Delay_LH_A1_S4 = $&delay_LH_A1_S4">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_HL_A1_S4 = $&delay_HL_A1_S4">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_A1_S4 = $&delay_A1_S4" >> "4_bit_Multiplier_Pre_Layout_pd.txt"
echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo "Delay_LH_A1_S5 = $&delay_LH_A1_S5">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_HL_A1_S5 = $&delay_HL_A1_S5">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_A1_S5 = $&delay_A1_S5" >> "4_bit_Multiplier_Pre_Layout_pd.txt"
echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo "Delay_LH_A1_S6 = $&delay_LH_A1_S6">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_HL_A1_S6 = $&delay_HL_A1_S6">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_A1_S6 = $&delay_A1_S6" >> "4_bit_Multiplier_Pre_Layout_pd.txt"
echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo "Delay_LH_A1_C = $&delay_LH_A1_C">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_HL_A1_C = $&delay_HL_A1_C">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_A1_C = $&delay_A1_C" >> "4_bit_Multiplier_Pre_Layout_pd.txt"
echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

****************************************************

* A2
meas tran delay_LH_A2_S0
+ TRIG v(A2) val = 0.5 rise = 3
+ TARG v(S0) val = 0.5 rise = 5
meas tran delay_HL_A2_S0
+ TRIG v(A2) val = 0.5 rise = 1
+ TARG v(S0) val = 0.5 fall = 2
let delay_A2_S0 = (delay_LH_A2_S0+delay_HL_A2_S0)/2

meas tran delay_LH_A2_S2
+ TRIG v(A2) val = 0.5 rise = 3
+ TARG v(S2) val = 0.5 rise = 6
meas tran delay_HL_A2_S2
+ TRIG v(A2) val = 0.5 rise = 2
+ TARG v(S2) val = 0.5 fall = 4
let delay_A2_S2 = (delay_LH_A2_S2+delay_HL_A2_S2)/2

meas tran delay_LH_A2_S3
+ TRIG v(A2) val = 0.5 rise = 2
+ TARG v(S3) val = 0.5 rise = 5
meas tran delay_HL_A2_S3
+ TRIG v(A2) val = 0.5 rise = 1
+ TARG v(S3) val = 0.5 fall = 1
let delay_A2_S3 = (delay_LH_A2_S3+delay_HL_A2_S3)/2

meas tran delay_LH_A2_S4
+ TRIG v(A2) val = 0.5 rise = 1
+ TARG v(S4) val = 0.5 rise = 1
meas tran delay_HL_A2_S4
+ TRIG v(A2) val = 0.5 rise = 3
+ TARG v(S4) val = 0.5 fall = 3
let delay_A2_S4 = (delay_LH_A2_S4+delay_HL_A2_S4)/2

meas tran delay_LH_A2_S5
+ TRIG v(A2) val = 0.5 fall = 2
+ TARG v(S5) val = 0.5 rise = 3
meas tran delay_HL_A2_S5
+ TRIG v(A2) val = 0.5 fall = 1
+ TARG v(S5) val = 0.5 fall = 2
let delay_A2_S5 = (delay_LH_A2_S5+delay_HL_A2_S5)/2

meas tran delay_LH_A2_S6
+ TRIG v(A2) val = 0.5 fall = 2
+ TARG v(S6) val = 0.5 rise = 3
meas tran delay_HL_A2_S6
+ TRIG v(A2) val = 0.5 rise = 1
+ TARG v(S6) val = 0.5 fall = 1
let delay_A2_S6 = (delay_LH_A2_S6+delay_HL_A2_S6)/2

meas tran delay_LH_A2_C
+ TRIG v(A2) val = 0.5 rise = 1
+ TARG v(C) val = 0.5 rise = 1
meas tran delay_HL_A2_C
+ TRIG v(A2) val = 0.5 fall = 1
+ TARG v(C) val = 0.5 fall = 1 
let delay_A2_C = (delay_LH_A2_C+delay_HL_A2_C)/2 

echo "A2">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo "Delay_LH_A2_S0 = $&delay_LH_A2_S0">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_HL_A2_S0 = $&delay_HL_A2_S0">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_A2_S0 = $&delay_A2_S0" >> "4_bit_Multiplier_Pre_Layout_pd.txt"
echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo "Delay_LH_A2_S2 = $&delay_LH_A2_S2">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_HL_A2_S2 = $&delay_HL_A2_S2">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_A2_S2 = $&delay_A2_S2" >> "4_bit_Multiplier_Pre_Layout_pd.txt"
echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo "Delay_LH_A2_S3 = $&delay_LH_A2_S3">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_HL_A2_S3 = $&delay_HL_A2_S3">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_A2_S3 = $&delay_A2_S3" >> "4_bit_Multiplier_Pre_Layout_pd.txt"
echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo "Delay_LH_A2_S4 = $&delay_LH_A2_S4">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_HL_A2_S4 = $&delay_HL_A2_S4">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_A2_S4 = $&delay_A2_S4" >> "4_bit_Multiplier_Pre_Layout_pd.txt"
echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo "Delay_LH_A2_S5 = $&delay_LH_A2_S5">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_HL_A2_S5 = $&delay_HL_A2_S5">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_A2_S5 = $&delay_A2_S5" >> "4_bit_Multiplier_Pre_Layout_pd.txt"
echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo "Delay_LH_A2_S6 = $&delay_LH_A2_S6">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_HL_A2_S6 = $&delay_HL_A2_S6">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_A2_S6 = $&delay_A2_S6" >> "4_bit_Multiplier_Pre_Layout_pd.txt"
echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo "Delay_LH_A2_C = $&delay_LH_A2_C">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_HL_A2_C = $&delay_HL_A2_C">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_A2_C = $&delay_A2_C" >> "4_bit_Multiplier_Pre_Layout_pd.txt"
echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

**************************************************

*A3
meas tran delay_LH_A3_S0
+ TRIG v(A3) val = 0.5 fall = 1
+ TARG v(S0) val = 0.5 fall = 4
meas tran delay_HL_A3_S0
+ TRIG v(A3) val = 0.5 rise = 1
+ TARG v(S0) val = 0.5 fall = 2
let delay_A3_S0 = (delay_LH_A3_S0+delay_HL_A3_S0)/2

meas tran delay_LH_A3_S2
+ TRIG v(A3) val = 0.5 rise = 2
+ TARG v(S2) val = 0.5 fall = 4
meas tran delay_HL_A3_S2
+ TRIG v(A3) val = 0.5 rise = 2
+ TARG v(S2) val = 0.5 fall = 4
let delay_A3_S2 = (delay_LH_A3_S2+delay_HL_A3_S2)/2

meas tran delay_LH_A3_S3
+ TRIG v(A3) val = 0.5 rise = 2
+ TARG v(S3) val = 0.5 rise = 5
meas tran delay_HL_A3_S3
+ TRIG v(A3) val = 0.5 rise = 1
+ TARG v(S3) val = 0.5 fall = 1
let delay_A3_S3 = (delay_LH_A3_S3+delay_HL_A3_S3)/2

meas tran delay_LH_A3_S4
+ TRIG v(A3) val = 0.5 rise = 1
+ TARG v(S4) val = 0.5 rise = 1
meas tran delay_HL_A3_S4
+ TRIG v(A3) val = 0.5 fall = 1
+ TARG v(S4) val = 0.5 fall = 2
let delay_A3_S4 = (delay_LH_A3_S4+delay_HL_A3_S4)/2

meas tran delay_LH_A3_S6
+ TRIG v(A3) val = 0.5 rise = 1
+ TARG v(S6) val = 0.5 rise = 1
meas tran delay_HL_A3_S6
+ TRIG v(A3) val = 0.5 fall = 1
+ TARG v(S6) val = 0.5 fall = 2
let delay_A3_S6 = (delay_LH_A3_S6+delay_HL_A3_S6)/2

meas tran delay_LH_A3_C
+ TRIG v(A3) val = 0.5 rise = 1
+ TARG v(C) val = 0.5 rise = 1
meas tran delay_HL_A3_C
+ TRIG v(A3) val = 0.5 fall = 1
+ TARG v(C) val = 0.5 fall = 1
let delay_A3_C = (delay_LH_A3_C+delay_HL_A3_C)/2 

echo "A3">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo "Delay_LH_A3_S0 = $&delay_LH_A3_S0">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_HL_A3_S0 = $&delay_HL_A3_S0">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_A3_S0 = $&delay_A3_S0" >> "4_bit_Multiplier_Pre_Layout_pd.txt"
echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo "Delay_LH_A3_S2 = $&delay_LH_A3_S2">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_HL_A3_S2 = $&delay_HL_A3_S2">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_A3_S2 = $&delay_A3_S2" >> "4_bit_Multiplier_Pre_Layout_pd.txt"
echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo "Delay_LH_A3_S3 = $&delay_LH_A3_S3">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_HL_A3_S3 = $&delay_HL_A3_S3">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_A3_S3 = $&delay_A3_S3" >> "4_bit_Multiplier_Pre_Layout_pd.txt"
echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo "Delay_LH_A3_S4 = $&delay_LH_A3_S4">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_HL_A3_S4 = $&delay_HL_A3_S4">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_A3_S4 = $&delay_A3_S4" >> "4_bit_Multiplier_Pre_Layout_pd.txt"
echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo "Delay_LH_A3_S6 = $&delay_LH_A3_S6">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_HL_A3_S6 = $&delay_HL_A3_S6">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_A3_S6 = $&delay_A3_S6" >> "4_bit_Multiplier_Pre_Layout_pd.txt"
echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo "Delay_LH_A3_C = $&delay_LH_A3_C">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_HL_A3_C = $&delay_HL_A3_C">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_A3_C = $&delay_A3_C" >> "4_bit_Multiplier_Pre_Layout_pd.txt"
echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

*****************************************************

*B0
meas tran delay_LH_B0_S0
+ TRIG v(B0) val = 0.5 rise = 1
+ TARG v(S0) val = 0.5 rise = 1
meas tran delay_HL_B0_S0
+ TRIG v(B0) val = 0.5 fall = 1
+ TARG v(S0) val = 0.5 fall = 1
let delay_B0_S0 = (delay_LH_B0_S0+delay_HL_B0_S0)/2

meas tran delay_LH_B0_S2
+ TRIG v(B0) val = 0.5 fall = 1
+ TARG v(S2) val = 0.5 rise = 1
meas tran delay_HL_B0_S2
+ TRIG v(B0) val = 0.5 rise = 2
+ TARG v(S2) val = 0.5 fall = 1
let delay_B0_S2 = (delay_LH_B0_S2+delay_HL_B0_S2)/2

meas tran delay_LH_B0_S3
+ TRIG v(B0) val = 0.5 fall = 4
+ TARG v(S3) val = 0.5 rise = 4
meas tran delay_HL_B0_S3
+ TRIG v(B0) val = 0.5 rise = 4
+ TARG v(S3) val = 0.5 fall = 3
let delay_B0_S3 = (delay_LH_B0_S3+delay_HL_B0_S3)/2

meas tran delay_LH_B0_S4
+ TRIG v(B0) val = 0.5 fall = 2
+ TARG v(S4) val = 0.5 rise = 1
meas tran delay_HL_B0_S4
+ TRIG v(B0) val = 0.5 rise = 3
+ TARG v(S4) val = 0.5 fall = 1
let delay_B0_S4 = (delay_LH_B0_S4+delay_HL_B0_S4)/2

meas tran delay_LH_B0_S5
+ TRIG v(B0) val = 0.5 fall = 6
+ TARG v(S5) val = 0.5 rise = 4
meas tran delay_HL_B0_S5
+ TRIG v(B0) val = 0.5 rise = 6
+ TARG v(S5) val = 0.5 fall = 3
let delay_B0_S5 = (delay_LH_B0_S5+delay_HL_B0_S5)/2

meas tran delay_LH_B0_S6
+ TRIG v(B0) val = 0.5 fall = 3
+ TARG v(S6) val = 0.5 rise = 2
meas tran delay_HL_B0_S6
+ TRIG v(B0) val = 0.5 rise = 6
+ TARG v(S6) val = 0.5 fall = 3
let delay_B0_S6 = (delay_LH_B0_S6+delay_HL_B0_S6)/2

meas tran delay_LH_B0_C
+ TRIG v(B0) val = 0.5 fall = 2
+ TARG v(C) val = 0.5 rise = 1
meas tran delay_HL_B0_C 
+ TRIG v(B0) val = 0.5 rise = 8
+ TARG v(C) val = 0.5 fall = 3 
let delay_B0_C = (delay_LH_B0_C+delay_HL_B0_C)/2 

echo "B0">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo "Delay_LH_B0_S0 = $&delay_LH_B0_S0">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_HL_B0_S0 = $&delay_HL_B0_S0">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_B0_S0 = $&delay_B0_S0" >> "4_bit_Multiplier_Pre_Layout_pd.txt"
echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo "Delay_LH_B0_S2 = $&delay_LH_B0_S2">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_HL_B0_S2 = $&delay_HL_B0_S2">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_B0_S2 = $&delay_B0_S2" >> "4_bit_Multiplier_Pre_Layout_pd.txt"
echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo "Delay_LH_B0_S3 = $&delay_LH_B0_S3">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_HL_B0_S3 = $&delay_HL_B0_S3">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_B0_S3 = $&delay_B0_S3" >> "4_bit_Multiplier_Pre_Layout_pd.txt"
echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo "Delay_LH_B0_S4 = $&delay_LH_B0_S4">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_HL_B0_S4 = $&delay_HL_B0_S4">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_B0_S4 = $&delay_B0_S4" >> "4_bit_Multiplier_Pre_Layout_pd.txt"
echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo "Delay_LH_B0_S5 = $&delay_LH_B0_S5">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_HL_B0_S5 = $&delay_HL_B0_S5">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_B0_S5 = $&delay_B0_S5" >> "4_bit_Multiplier_Pre_Layout_pd.txt"
echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo "Delay_LH_B0_S6 = $&delay_LH_B0_S6">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_HL_B0_S6 = $&delay_HL_B0_S6">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_B0_S6 = $&delay_B0_S6" >> "4_bit_Multiplier_Pre_Layout_pd.txt"
echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo "Delay_LH_B0_C = $&delay_LH_B0_C">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_HL_B0_C = $&delay_HL_B0_C">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_B0_C = $&delay_B0_C" >> "4_bit_Multiplier_Pre_Layout_pd.txt"
echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

*************************************************

*B1
meas tran delay_LH_B1_S0
+ TRIG v(B1) val = 0.5 fall = 3
+ TARG v(S0) val = 0.5 rise = 6
meas tran delay_HL_B1_S0
+ TRIG v(B1) val = 0.5 rise = 1
+ TARG v(S0) val = 0.5 fall = 1
let delay_B1_S0 = (delay_LH_B1_S0+delay_HL_B1_S0)/2

meas tran delay_LH_B1_S2
+ TRIG v(B1) val = 0.5 fall = 2
+ TARG v(S2) val = 0.5 rise = 5
meas tran delay_HL_B1_S2
+ TRIG v(B1) val = 0.5 rise = 3
+ TARG v(S2) val = 0.5 fall = 7
let delay_B1_S2 = (delay_LH_B1_S2+delay_HL_B1_S2)/2

meas tran delay_LH_B1_S3 
+ TRIG v(B1) val = 0.5 fall = 2
+ TARG v(S3) val = 0.5 rise = 5
meas tran delay_HL_B1_S3
+ TRIG v(B1) val = 0.5 rise = 2
+ TARG v(S3) val = 0.5 fall = 2
let delay_B1_S3 = (delay_LH_B1_S3+delay_HL_B1_S3)/2

meas tran delay_LH_B1_S4
+ TRIG v(B1) val = 0.5 fall = 1
+ TARG v(S4) val = 0.5 rise = 1
meas tran delay_HL_B1_S4
+ TRIG v(B1) val = 0.5 rise = 3
+ TARG v(S4) val = 0.5 fall = 4
let delay_B1_S4 = (delay_LH_B1_S4+delay_HL_B1_S4)/2

meas tran delay_LH_B1_S5 
+ TRIG v(B1) val = 0.5 fall = 3
+ TARG v(S5) val = 0.5 rise = 5
meas tran delay_HL_B1_S5
+ TRIG v(B1) val = 0.5 rise = 2
+ TARG v(S5) val = 0.5 fall = 1
let delay_B1_S5 = (delay_LH_B1_S5+delay_HL_B1_S5)/2

meas tran delay_LH_B1_S6
+ TRIG v(B1) val = 0.5 fall = 1
+ TARG v(S6) val = 0.5 rise = 1
meas tran delay_HL_B1_S6
+ TRIG v(B1) val = 0.5 rise = 4
+ TARG v(S6) val = 0.5 fall = 6
let delay_B1_S6 = (delay_LH_B1_S6+delay_HL_B1_S6)/2

meas tran delay_LH_B1_C
+ TRIG v(B1) val = 0.5 fall = 1
+ TARG v(C) val = 0.5 rise = 1
meas tran delay_HL_B1_C 
+ TRIG v(B1) val = 0.5 rise = 4
+ TARG v(C) val = 0.5 rise = 3 
let delay_B1_C = (delay_LH_B1_C+delay_HL_B1_C)/2 

echo "B1">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo "Delay_LH_B1_S0 = $&delay_LH_B1_S0">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_HL_B1_S0 = $&delay_HL_B1_S0">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_B1_S0 = $&delay_B1_S0" >> "4_bit_Multiplier_Pre_Layout_pd.txt"
echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo "Delay_LH_B1_S2 = $&delay_LH_B1_S2">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_HL_B1_S2 = $&delay_HL_B1_S2">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_B1_S2 = $&delay_B1_S2" >> "4_bit_Multiplier_Pre_Layout_pd.txt"
echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo "Delay_LH_B1_S3 = $&delay_LH_B1_S3">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_HL_B1_S3 = $&delay_HL_B1_S3">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_B1_S3 = $&delay_B1_S3" >> "4_bit_Multiplier_Pre_Layout_pd.txt"
echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo "Delay_LH_B1_S4 = $&delay_LH_B1_S4">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_HL_B1_S4 = $&delay_HL_B1_S4">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_B1_S4 = $&delay_B1_S4" >> "4_bit_Multiplier_Pre_Layout_pd.txt"
echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo "Delay_LH_B1_S5 = $&delay_LH_B1_S5">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_HL_B1_S5 = $&delay_HL_B1_S5">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_B1_S5 = $&delay_B1_S5" >> "4_bit_Multiplier_Pre_Layout_pd.txt"
echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo "Delay_LH_B1_S6 = $&delay_LH_B1_S6">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_HL_B1_S6 = $&delay_HL_B1_S6">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_B1_S6 = $&delay_B1_S6" >> "4_bit_Multiplier_Pre_Layout_pd.txt"
echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo "Delay_LH_B1_C = $&delay_LH_B1_C">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_HL_B1_C = $&delay_HL_B1_C">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_B1_C = $&delay_B1_C" >> "4_bit_Multiplier_Pre_Layout_pd.txt"
echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

**************************************************

*B2
meas tran delay_LH_B2_S0
+ TRIG v(B2) val = 0.5 rise = 1
+ TARG v(S0) val = 0.5 fall = 2
meas tran delay_HL_B2_S0
+ TRIG v(B2) val = 0.5 rise = 1
+ TARG v(S0) val = 0.5 fall = 2
let delay_B2_S0 = (delay_LH_B2_S0+delay_HL_B2_S0)/2

meas tran delay_LH_B2_S2
+ TRIG v(B2) val = 0.5 fall = 2
+ TARG v(S2) val = 0.5 rise = 8
meas tran delay_HL_B2_S2
+ TRIG v(B2) val = 0.5 fall = 1
+ TARG v(S2) val = 0.5 fall = 4
let delay_B2_S2 = (delay_LH_B2_S2+delay_HL_B2_S2)/2

meas tran delay_LH_B2_S3
+ TRIG v(B2) val = 0.5 fall = 1
+ TARG v(S3) val = 0.5 rise = 5
meas tran delay_HL_B2_S3
+ TRIG v(B2) val = 0.5 rise = 1
+ TARG v(S3) val = 0.5 fall = 1
let delay_B2_S3 = (delay_LH_B2_S3+delay_HL_B2_S3)/2

meas tran delay_LH_B2_S4
+ TRIG v(B2) val = 0.5 rise = 1
+ TARG v(S4) val = 0.5 rise = 1
meas tran delay_HL_B2_S4
+ TRIG v(B2) val = 0.5 fall = 2
+ TARG v(S4) val = 0.5 fall = 5
let delay_B2_S4 = (delay_LH_B2_S4+delay_HL_B2_S4)/2

meas tran delay_LH_B2_S5
+ TRIG v(B2) val = 0.5 rise = 2
+ TARG v(S5) val = 0.5 rise = 3
meas tran delay_HL_B2_S5
+ TRIG v(B2) val = 0.5 rise = 2
+ TARG v(S5) val = 0.5 rise = 3
let delay_B2_S5 = (delay_LH_B2_S5+delay_HL_B2_S5)/2

meas tran delay_LH_B2_S6
+ TRIG v(B2) val = 0.5 rise = 2
+ TARG v(S6) val = 0.5 rise = 3
meas tran delay_HL_B2_S6
+ TRIG v(B2) val = 0.5 rise = 1
+ TARG v(S6) val = 0.5 fall = 1
let delay_B2_S6 = (delay_LH_B2_S6+delay_HL_B2_S6)/2

meas tran delay_LH_B2_C
+ TRIG v(B2) val = 0.5 rise = 1
+ TARG v(C) val = 0.5 rise = 1
meas tran delay_HL_B2_C
+ TRIG v(B2) val = 0.5 fall = 2
+ TARG v(C) val = 0.5 fall = 2 
let delay_B2_C = (delay_LH_B2_C+delay_HL_B2_C)/2 

echo "B2">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo "Delay_LH_B2_S0 = $&delay_LH_B2_S0">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_HL_B2_S0 = $&delay_HL_B2_S0">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_B2_S0 = $&delay_B2_S0" >> "4_bit_Multiplier_Pre_Layout_pd.txt"
echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo "Delay_LH_B2_S2 = $&delay_LH_B2_S2">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_HL_B2_S2 = $&delay_HL_B2_S2">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_B2_S2 = $&delay_B2_S2" >> "4_bit_Multiplier_Pre_Layout_pd.txt"
echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo "Delay_LH_B2_S3 = $&delay_LH_B2_S3">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_HL_B2_S3 = $&delay_HL_B2_S3">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_B2_S3 = $&delay_B2_S3" >> "4_bit_Multiplier_Pre_Layout_pd.txt"
echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo "Delay_LH_B2_S4 = $&delay_LH_B2_S4">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_HL_B2_S4 = $&delay_HL_B2_S4">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_B2_S4 = $&delay_B2_S4" >> "4_bit_Multiplier_Pre_Layout_pd.txt"
echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo "Delay_LH_B2_S5 = $&delay_LH_B2_S5">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_HL_B2_S5 = $&delay_HL_B2_S5">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_B2_S5 = $&delay_B2_S5" >> "4_bit_Multiplier_Pre_Layout_pd.txt"
echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo "Delay_LH_B2_S6 = $&delay_LH_B2_S6">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_HL_B2_S6 = $&delay_HL_B2_S6">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_B2_S6 = $&delay_B2_S6" >> "4_bit_Multiplier_Pre_Layout_pd.txt"
echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo "Delay_LH_B2_C = $&delay_LH_B2_C">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_HL_B2_C = $&delay_HL_B2_C">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_B2_C = $&delay_B2_C" >> "4_bit_Multiplier_Pre_Layout_pd.txt"
echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

**************************************************

*B3
meas tran delay_LH_B3_S0
+ TRIG v(B3) val = 0.5 rise = 1
+ TARG v(S0) val = 0.5 fall = 2
meas tran delay_HL_B3_S0
+ TRIG v(B3) val = 0.5 fall = 2
+ TARG v(S0) val = 0.5 rise = 5
let delay_B3_S0 = (delay_LH_B3_S0+delay_HL_B3_S0)/2

meas tran delay_LH_B3_S2
+ TRIG v(B3) val = 0.5 fall = 3
+ TARG v(S2) val = 0.5 rise = 8
meas tran delay_HL_B3_S2
+ TRIG v(B3) val = 0.5 fall = 1
+ TARG v(S2) val = 0.5 fall = 4
let delay_B3_S2 = (delay_LH_B3_S2+delay_HL_B3_S2)/2

meas tran delay_LH_B3_S3
+ TRIG v(B3) val = 0.5 rise = 3
+ TARG v(S3) val = 0.5 rise = 6
meas tran delay_HL_B3_S3
+ TRIG v(B3) val = 0.5 rise = 1
+ TARG v(S3) val = 0.5 fall = 1
let delay_B3_S3 = (delay_LH_B3_S3+delay_HL_B3_S3)/2

meas tran delay_LH_B3_S4
+ TRIG v(B3) val = 0.5 fall = 3
+ TARG v(S4) val = 0.5 rise = 6
meas tran delay_HL_B3_S4
+ TRIG v(B3) val = 0.5 fall = 2
+ TARG v(S4) val = 0.5 fall = 3
let delay_B3_S4 = (delay_LH_B3_S4+delay_HL_B3_S4)/2

meas tran delay_LH_B3_S5
+ TRIG v(B3) val = 0.5 rise = 2
+ TARG v(S5) val = 0.5 rise = 3
meas tran delay_HL_B3_S5
+ TRIG v(B3) val = 0.5 fall = 2
+ TARG v(S5) val = 0.5 fall = 3
let delay_B3_S5 = (delay_LH_B3_S5+delay_HL_B3_S5)/2

meas tran delay_LH_B3_S6
+ TRIG v(B3) val = 0.5 rise = 1
+ TARG v(S6) val = 0.5 rise = 1
meas tran delay_HL_B3_S6
+ TRIG v(B3) val = 0.5 rise = 3
+ TARG v(S6) val = 0.5 fall = 4
let delay_B3_S6 = (delay_LH_B3_S6+delay_HL_B3_S6)/2

meas tran delay_LH_B3_C
+ TRIG v(B3) val = 0.5 rise = 1
+ TARG v(C) val = 0.5 rise = 1
meas tran delay_HL_B3_C
+ TRIG v(B3) val = 0.5 rise = 3
+ TARG v(C) val = 0.5 rise = 2 
let delay_B3_C = (delay_LH_B3_C+delay_HL_B3_C)/2 

echo "B3">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo "Delay_LH_B3_S0 = $&delay_LH_B3_S0">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_HL_B3_S0 = $&delay_HL_B3_S0">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_B3_S0 = $&delay_B3_S0" >> "4_bit_Multiplier_Pre_Layout_pd.txt"
echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo "Delay_LH_B3_S2 = $&delay_LH_B3_S2">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_HL_B3_S2 = $&delay_HL_B3_S2">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_B3_S2 = $&delay_B3_S2" >> "4_bit_Multiplier_Pre_Layout_pd.txt"
echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo "Delay_LH_B3_S3 = $&delay_LH_B3_S3">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_HL_B3_S3 = $&delay_HL_B3_S3">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_B3_S3 = $&delay_B3_S3" >> "4_bit_Multiplier_Pre_Layout_pd.txt"
echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo "Delay_LH_B3_S4 = $&delay_LH_B3_S4">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_HL_B3_S4 = $&delay_HL_B3_S4">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_B3_S4 = $&delay_B3_S4" >> "4_bit_Multiplier_Pre_Layout_pd.txt"
echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo "Delay_LH_B3_S5 = $&delay_LH_B3_S5">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_HL_B3_S5 = $&delay_HL_B3_S5">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_B3_S5 = $&delay_B3_S5" >> "4_bit_Multiplier_Pre_Layout_pd.txt"
echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo "Delay_LH_B3_S6 = $&delay_LH_B3_S6">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_HL_B3_S6 = $&delay_HL_B3_S6">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_B3_S6 = $&delay_B3_S6" >> "4_bit_Multiplier_Pre_Layout_pd.txt"
echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo "Delay_LH_B3_C = $&delay_LH_B3_C">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_HL_B3_C = $&delay_HL_B3_C">>"4_bit_Multiplier_Pre_Layout_pd.txt"
echo "Delay_B3_C = $&delay_B3_C" >> "4_bit_Multiplier_Pre_Layout_pd.txt"
echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

echo " ">>"4_bit_Multiplier_Pre_Layout_pd.txt"

****************************************************
hardcopy 4_Bit_Multiplier_Pre_Layout_A.eps V(A0)+6 V(A1)+4 V(A2)+2 V(A3)
hardcopy 4_Bit_Multiplier_Pre_Layout_B.eps V(B0)+6 V(B1)+4 V(B2)+2 V(B3)
hardcopy 4_Bit_Multiplier_Pre_Layout_OUT.eps V(C)+16 V(S6)+14 V(S5)+12 V(S4)+10 V(S3)+8 V(S2)+6 V(S1)+4 V(S0)+2

.endc