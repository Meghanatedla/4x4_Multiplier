magic
tech scmos
timestamp 1667670020
<< nwell >>
rect -88 -472 58 -437
<< ntransistor >>
rect -77 -513 -75 -509
rect -69 -513 -67 -509
rect -63 -513 -61 -509
rect -55 -513 -53 -509
rect -47 -513 -45 -509
rect -39 -513 -37 -509
rect -33 -513 -31 -509
rect -27 -513 -25 -509
rect -16 -513 -14 -509
rect -3 -513 -1 -509
rect 5 -513 7 -509
rect 13 -513 15 -509
rect 25 -513 27 -509
rect 44 -513 46 -509
rect -74 -522 -70 -520
<< ptransistor >>
rect -77 -466 -75 -458
rect -69 -466 -67 -458
rect -63 -466 -61 -458
rect -55 -466 -53 -458
rect -47 -466 -45 -458
rect -39 -466 -37 -458
rect -33 -466 -31 -458
rect -27 -466 -25 -458
rect -16 -466 -14 -458
rect -3 -466 -1 -458
rect 5 -466 7 -458
rect 13 -466 15 -458
rect 25 -466 27 -458
rect 44 -466 46 -458
<< ndiffusion >>
rect -24 -509 -20 -497
rect -10 -509 -6 -497
rect -78 -513 -77 -509
rect -75 -513 -69 -509
rect -67 -513 -63 -509
rect -61 -513 -60 -509
rect -56 -513 -55 -509
rect -53 -513 -52 -509
rect -48 -513 -47 -509
rect -45 -513 -44 -509
rect -40 -513 -39 -509
rect -37 -513 -33 -509
rect -31 -513 -27 -509
rect -25 -513 -16 -509
rect -14 -513 -3 -509
rect -1 -513 0 -509
rect 4 -513 5 -509
rect 7 -513 8 -509
rect 12 -513 13 -509
rect 15 -513 18 -509
rect 22 -513 25 -509
rect 27 -513 30 -509
rect 43 -513 44 -509
rect 46 -513 47 -509
rect -74 -520 -70 -513
rect -74 -526 -70 -522
<< pdiffusion >>
rect -74 -458 -70 -447
rect -78 -466 -77 -458
rect -75 -466 -69 -458
rect -67 -466 -63 -458
rect -61 -466 -60 -458
rect -56 -466 -55 -458
rect -53 -466 -52 -458
rect -48 -466 -47 -458
rect -45 -466 -44 -458
rect -40 -466 -39 -458
rect -37 -466 -33 -458
rect -31 -466 -27 -458
rect -25 -466 -24 -458
rect -20 -466 -16 -458
rect -14 -466 -10 -458
rect -6 -466 -3 -458
rect -1 -466 0 -458
rect 4 -466 5 -458
rect 7 -466 8 -458
rect 12 -466 13 -458
rect 15 -466 18 -458
rect 22 -466 25 -458
rect 27 -466 30 -458
rect 43 -466 44 -458
rect 46 -466 47 -458
rect 51 -466 52 -458
<< ndcontact >>
rect -24 -497 -20 -493
rect -10 -497 -6 -493
rect -82 -513 -78 -509
rect -60 -513 -56 -509
rect -52 -513 -48 -509
rect -44 -513 -40 -509
rect 0 -513 4 -509
rect 8 -513 12 -509
rect 18 -513 22 -509
rect 30 -513 34 -509
rect 39 -513 43 -509
rect 47 -513 51 -509
rect -74 -530 -70 -526
<< pdcontact >>
rect -74 -447 -70 -443
rect -82 -466 -78 -458
rect -60 -466 -56 -458
rect -52 -466 -48 -458
rect -44 -466 -40 -458
rect -24 -466 -20 -458
rect -10 -466 -6 -458
rect 0 -466 4 -458
rect 8 -466 12 -458
rect 18 -466 22 -458
rect 30 -466 34 -458
rect 39 -466 43 -458
rect 47 -466 51 -458
<< polysilicon >>
rect -47 -445 -45 -435
rect -77 -458 -75 -455
rect -69 -447 7 -445
rect -69 -458 -67 -447
rect -63 -452 -45 -450
rect -63 -458 -61 -452
rect -55 -458 -53 -455
rect -47 -458 -45 -452
rect -39 -458 -37 -455
rect -33 -458 -31 -447
rect -27 -458 -25 -455
rect -16 -458 -14 -455
rect -3 -458 -1 -455
rect 5 -458 7 -447
rect 13 -458 15 -455
rect 25 -458 27 -454
rect 44 -458 46 -455
rect -77 -468 -75 -466
rect -69 -468 -67 -466
rect -77 -470 -67 -468
rect -77 -509 -75 -470
rect -69 -509 -67 -470
rect -63 -509 -61 -466
rect -55 -509 -53 -466
rect -47 -468 -45 -466
rect -39 -468 -37 -466
rect -47 -470 -37 -468
rect -47 -492 -45 -470
rect -47 -509 -45 -497
rect -39 -509 -37 -470
rect -33 -509 -31 -466
rect -27 -509 -25 -466
rect -16 -501 -14 -466
rect -16 -509 -14 -506
rect -3 -509 -1 -466
rect 5 -509 7 -466
rect 13 -509 15 -466
rect 25 -509 27 -466
rect 44 -509 46 -466
rect -86 -520 -84 -514
rect -77 -516 -75 -513
rect -69 -516 -67 -513
rect -63 -516 -61 -513
rect -55 -520 -53 -513
rect -47 -516 -45 -513
rect -39 -516 -37 -513
rect -33 -516 -31 -513
rect -27 -520 -25 -513
rect -16 -516 -14 -513
rect -3 -520 -1 -513
rect 5 -516 7 -513
rect 13 -516 15 -513
rect 25 -516 27 -513
rect 44 -516 46 -513
rect -86 -522 -74 -520
rect -70 -522 -1 -520
<< polycontact >>
rect -48 -497 -43 -492
rect -16 -506 -11 -501
rect 21 -486 25 -482
rect 15 -497 20 -492
rect 39 -505 44 -500
<< metal1 >>
rect -88 -447 -74 -443
rect -70 -447 58 -443
rect -82 -454 -48 -450
rect -82 -458 -78 -454
rect -52 -458 -48 -454
rect -44 -458 -40 -447
rect 0 -458 4 -447
rect 18 -458 22 -447
rect 39 -458 43 -447
rect -60 -501 -56 -466
rect -24 -482 -20 -466
rect -10 -469 -6 -466
rect 8 -469 12 -466
rect -10 -473 12 -469
rect 30 -478 34 -466
rect -24 -486 21 -482
rect -24 -493 -20 -486
rect -6 -497 12 -493
rect -60 -505 -16 -501
rect -60 -509 -56 -505
rect 8 -509 12 -497
rect 30 -509 34 -483
rect 47 -490 51 -466
rect 60 -482 64 -478
rect 47 -494 64 -490
rect 47 -509 51 -494
rect -82 -518 -78 -513
rect -52 -518 -48 -513
rect -82 -522 -48 -518
rect -44 -526 -40 -513
rect 0 -526 4 -513
rect 18 -526 22 -513
rect 39 -526 43 -513
rect -87 -530 -74 -526
rect -70 -530 51 -526
<< m2contact >>
rect 30 -483 35 -478
rect 55 -483 60 -478
<< pm12contact >>
rect -48 -497 -43 -492
rect 15 -497 20 -492
rect -16 -506 -11 -501
rect 39 -505 44 -500
<< metal2 >>
rect -24 -493 -20 -435
rect 35 -482 55 -478
rect -43 -497 15 -493
rect -11 -505 39 -501
<< labels >>
rlabel metal1 -88 -447 -77 -443 1 VDD
rlabel metal1 -87 -530 -74 -526 1 GND
rlabel polysilicon -86 -516 -84 -514 1 C
rlabel polysilicon -47 -437 -45 -435 1 A
rlabel metal2 -24 -437 -20 -435 1 B
rlabel metal1 60 -482 64 -478 7 SUM
rlabel metal1 60 -494 64 -490 7 CARRY
<< end >>
