magic
tech scmos
timestamp 1669640817
<< nwell >>
rect -340 -3 -290 17
rect -219 -3 -169 17
rect -105 -3 -55 17
rect -5 -3 45 17
rect -440 -221 -390 -201
rect -282 -221 -232 -201
rect -143 -221 -93 -201
rect -25 -221 25 -201
rect -718 -389 -668 -369
rect -604 -395 -458 -360
rect -352 -395 -206 -360
rect -12 -389 38 -369
rect -775 -469 -751 -449
rect -733 -469 -677 -449
rect -69 -469 -45 -449
rect -27 -469 29 -449
rect -775 -521 -751 -501
rect -69 -521 -45 -501
rect -725 -707 -675 -687
rect -547 -707 -497 -687
rect -367 -707 -317 -687
rect -156 -707 -106 -687
rect -826 -865 -680 -830
rect -600 -865 -454 -830
rect -382 -865 -236 -830
rect 7 -859 57 -839
rect -50 -939 -26 -919
rect -8 -939 48 -919
rect -50 -991 -26 -971
rect -725 -1212 -675 -1192
rect -547 -1212 -497 -1192
rect -367 -1212 -317 -1192
rect -156 -1212 -106 -1192
rect -871 -1430 -725 -1395
rect -645 -1430 -499 -1395
rect -427 -1430 -281 -1395
rect 7 -1423 57 -1403
rect -50 -1503 -26 -1483
rect -8 -1503 48 -1483
rect -50 -1555 -26 -1535
<< ntransistor >>
rect -303 -16 -301 -12
rect -329 -25 -327 -21
rect -319 -25 -317 -21
rect -182 -16 -180 -12
rect -208 -25 -206 -21
rect -198 -25 -196 -21
rect -68 -16 -66 -12
rect -94 -25 -92 -21
rect -84 -25 -82 -21
rect 32 -16 34 -12
rect 6 -25 8 -21
rect 16 -25 18 -21
rect -403 -234 -401 -230
rect -429 -243 -427 -239
rect -419 -243 -417 -239
rect -245 -234 -243 -230
rect -271 -243 -269 -239
rect -261 -243 -259 -239
rect -106 -234 -104 -230
rect -132 -243 -130 -239
rect -122 -243 -120 -239
rect 12 -234 14 -230
rect -14 -243 -12 -239
rect -4 -243 -2 -239
rect -681 -402 -679 -398
rect -707 -411 -705 -407
rect -697 -411 -695 -407
rect 25 -402 27 -398
rect -1 -411 1 -407
rect 9 -411 11 -407
rect -593 -436 -591 -432
rect -585 -436 -583 -432
rect -579 -436 -577 -432
rect -571 -436 -569 -432
rect -563 -436 -561 -432
rect -555 -436 -553 -432
rect -549 -436 -547 -432
rect -543 -436 -541 -432
rect -532 -436 -530 -432
rect -519 -436 -517 -432
rect -511 -436 -509 -432
rect -503 -436 -501 -432
rect -491 -436 -489 -432
rect -472 -436 -470 -432
rect -341 -436 -339 -432
rect -333 -436 -331 -432
rect -327 -436 -325 -432
rect -319 -436 -317 -432
rect -311 -436 -309 -432
rect -303 -436 -301 -432
rect -297 -436 -295 -432
rect -291 -436 -289 -432
rect -280 -436 -278 -432
rect -267 -436 -265 -432
rect -259 -436 -257 -432
rect -251 -436 -249 -432
rect -239 -436 -237 -432
rect -220 -436 -218 -432
rect -590 -445 -586 -443
rect -338 -445 -334 -443
rect -764 -481 -762 -477
rect -58 -481 -56 -477
rect -764 -533 -762 -529
rect -720 -533 -718 -529
rect -711 -533 -709 -529
rect -702 -533 -700 -529
rect -692 -533 -690 -529
rect -58 -533 -56 -529
rect -14 -533 -12 -529
rect -5 -533 -3 -529
rect 4 -533 6 -529
rect 14 -533 16 -529
rect -688 -720 -686 -716
rect -714 -729 -712 -725
rect -704 -729 -702 -725
rect -510 -720 -508 -716
rect -536 -729 -534 -725
rect -526 -729 -524 -725
rect -330 -720 -328 -716
rect -356 -729 -354 -725
rect -346 -729 -344 -725
rect -119 -720 -117 -716
rect -145 -729 -143 -725
rect -135 -729 -133 -725
rect 44 -872 46 -868
rect 18 -881 20 -877
rect 28 -881 30 -877
rect -815 -906 -813 -902
rect -807 -906 -805 -902
rect -801 -906 -799 -902
rect -793 -906 -791 -902
rect -785 -906 -783 -902
rect -777 -906 -775 -902
rect -771 -906 -769 -902
rect -765 -906 -763 -902
rect -754 -906 -752 -902
rect -741 -906 -739 -902
rect -733 -906 -731 -902
rect -725 -906 -723 -902
rect -713 -906 -711 -902
rect -694 -906 -692 -902
rect -589 -906 -587 -902
rect -581 -906 -579 -902
rect -575 -906 -573 -902
rect -567 -906 -565 -902
rect -559 -906 -557 -902
rect -551 -906 -549 -902
rect -545 -906 -543 -902
rect -539 -906 -537 -902
rect -528 -906 -526 -902
rect -515 -906 -513 -902
rect -507 -906 -505 -902
rect -499 -906 -497 -902
rect -487 -906 -485 -902
rect -468 -906 -466 -902
rect -371 -906 -369 -902
rect -363 -906 -361 -902
rect -357 -906 -355 -902
rect -349 -906 -347 -902
rect -341 -906 -339 -902
rect -333 -906 -331 -902
rect -327 -906 -325 -902
rect -321 -906 -319 -902
rect -310 -906 -308 -902
rect -297 -906 -295 -902
rect -289 -906 -287 -902
rect -281 -906 -279 -902
rect -269 -906 -267 -902
rect -250 -906 -248 -902
rect -812 -915 -808 -913
rect -586 -915 -582 -913
rect -368 -915 -364 -913
rect -39 -951 -37 -947
rect -39 -1003 -37 -999
rect 5 -1003 7 -999
rect 14 -1003 16 -999
rect 23 -1003 25 -999
rect 33 -1003 35 -999
rect -688 -1225 -686 -1221
rect -714 -1234 -712 -1230
rect -704 -1234 -702 -1230
rect -510 -1225 -508 -1221
rect -536 -1234 -534 -1230
rect -526 -1234 -524 -1230
rect -330 -1225 -328 -1221
rect -356 -1234 -354 -1230
rect -346 -1234 -344 -1230
rect -119 -1225 -117 -1221
rect -145 -1234 -143 -1230
rect -135 -1234 -133 -1230
rect 44 -1436 46 -1432
rect 18 -1445 20 -1441
rect 28 -1445 30 -1441
rect -860 -1471 -858 -1467
rect -852 -1471 -850 -1467
rect -846 -1471 -844 -1467
rect -838 -1471 -836 -1467
rect -830 -1471 -828 -1467
rect -822 -1471 -820 -1467
rect -816 -1471 -814 -1467
rect -810 -1471 -808 -1467
rect -799 -1471 -797 -1467
rect -786 -1471 -784 -1467
rect -778 -1471 -776 -1467
rect -770 -1471 -768 -1467
rect -758 -1471 -756 -1467
rect -739 -1471 -737 -1467
rect -634 -1471 -632 -1467
rect -626 -1471 -624 -1467
rect -620 -1471 -618 -1467
rect -612 -1471 -610 -1467
rect -604 -1471 -602 -1467
rect -596 -1471 -594 -1467
rect -590 -1471 -588 -1467
rect -584 -1471 -582 -1467
rect -573 -1471 -571 -1467
rect -560 -1471 -558 -1467
rect -552 -1471 -550 -1467
rect -544 -1471 -542 -1467
rect -532 -1471 -530 -1467
rect -513 -1471 -511 -1467
rect -416 -1471 -414 -1467
rect -408 -1471 -406 -1467
rect -402 -1471 -400 -1467
rect -394 -1471 -392 -1467
rect -386 -1471 -384 -1467
rect -378 -1471 -376 -1467
rect -372 -1471 -370 -1467
rect -366 -1471 -364 -1467
rect -355 -1471 -353 -1467
rect -342 -1471 -340 -1467
rect -334 -1471 -332 -1467
rect -326 -1471 -324 -1467
rect -314 -1471 -312 -1467
rect -295 -1471 -293 -1467
rect -857 -1480 -853 -1478
rect -631 -1480 -627 -1478
rect -413 -1480 -409 -1478
rect -39 -1515 -37 -1511
rect -39 -1567 -37 -1563
rect 5 -1567 7 -1563
rect 14 -1567 16 -1563
rect 23 -1567 25 -1563
rect 33 -1567 35 -1563
<< ptransistor >>
rect -329 3 -327 11
rect -319 3 -317 11
rect -303 3 -301 11
rect -208 3 -206 11
rect -198 3 -196 11
rect -182 3 -180 11
rect -94 3 -92 11
rect -84 3 -82 11
rect -68 3 -66 11
rect 6 3 8 11
rect 16 3 18 11
rect 32 3 34 11
rect -429 -215 -427 -207
rect -419 -215 -417 -207
rect -403 -215 -401 -207
rect -271 -215 -269 -207
rect -261 -215 -259 -207
rect -245 -215 -243 -207
rect -132 -215 -130 -207
rect -122 -215 -120 -207
rect -106 -215 -104 -207
rect -14 -215 -12 -207
rect -4 -215 -2 -207
rect 12 -215 14 -207
rect -707 -383 -705 -375
rect -697 -383 -695 -375
rect -681 -383 -679 -375
rect -593 -389 -591 -381
rect -585 -389 -583 -381
rect -579 -389 -577 -381
rect -571 -389 -569 -381
rect -563 -389 -561 -381
rect -555 -389 -553 -381
rect -549 -389 -547 -381
rect -543 -389 -541 -381
rect -532 -389 -530 -381
rect -519 -389 -517 -381
rect -511 -389 -509 -381
rect -503 -389 -501 -381
rect -491 -389 -489 -381
rect -472 -389 -470 -381
rect -341 -389 -339 -381
rect -333 -389 -331 -381
rect -327 -389 -325 -381
rect -319 -389 -317 -381
rect -311 -389 -309 -381
rect -303 -389 -301 -381
rect -297 -389 -295 -381
rect -291 -389 -289 -381
rect -280 -389 -278 -381
rect -267 -389 -265 -381
rect -259 -389 -257 -381
rect -251 -389 -249 -381
rect -239 -389 -237 -381
rect -220 -389 -218 -381
rect -1 -383 1 -375
rect 9 -383 11 -375
rect 25 -383 27 -375
rect -764 -463 -762 -455
rect -721 -463 -719 -455
rect -711 -463 -709 -455
rect -701 -463 -699 -455
rect -692 -463 -690 -455
rect -764 -515 -762 -507
rect -58 -463 -56 -455
rect -15 -463 -13 -455
rect -5 -463 -3 -455
rect 5 -463 7 -455
rect 14 -463 16 -455
rect -58 -515 -56 -507
rect -714 -701 -712 -693
rect -704 -701 -702 -693
rect -688 -701 -686 -693
rect -536 -701 -534 -693
rect -526 -701 -524 -693
rect -510 -701 -508 -693
rect -356 -701 -354 -693
rect -346 -701 -344 -693
rect -330 -701 -328 -693
rect -145 -701 -143 -693
rect -135 -701 -133 -693
rect -119 -701 -117 -693
rect -815 -859 -813 -851
rect -807 -859 -805 -851
rect -801 -859 -799 -851
rect -793 -859 -791 -851
rect -785 -859 -783 -851
rect -777 -859 -775 -851
rect -771 -859 -769 -851
rect -765 -859 -763 -851
rect -754 -859 -752 -851
rect -741 -859 -739 -851
rect -733 -859 -731 -851
rect -725 -859 -723 -851
rect -713 -859 -711 -851
rect -694 -859 -692 -851
rect -589 -859 -587 -851
rect -581 -859 -579 -851
rect -575 -859 -573 -851
rect -567 -859 -565 -851
rect -559 -859 -557 -851
rect -551 -859 -549 -851
rect -545 -859 -543 -851
rect -539 -859 -537 -851
rect -528 -859 -526 -851
rect -515 -859 -513 -851
rect -507 -859 -505 -851
rect -499 -859 -497 -851
rect -487 -859 -485 -851
rect -468 -859 -466 -851
rect -371 -859 -369 -851
rect -363 -859 -361 -851
rect -357 -859 -355 -851
rect -349 -859 -347 -851
rect -341 -859 -339 -851
rect -333 -859 -331 -851
rect -327 -859 -325 -851
rect -321 -859 -319 -851
rect -310 -859 -308 -851
rect -297 -859 -295 -851
rect -289 -859 -287 -851
rect -281 -859 -279 -851
rect -269 -859 -267 -851
rect -250 -859 -248 -851
rect 18 -853 20 -845
rect 28 -853 30 -845
rect 44 -853 46 -845
rect -39 -933 -37 -925
rect 4 -933 6 -925
rect 14 -933 16 -925
rect 24 -933 26 -925
rect 33 -933 35 -925
rect -39 -985 -37 -977
rect -714 -1206 -712 -1198
rect -704 -1206 -702 -1198
rect -688 -1206 -686 -1198
rect -536 -1206 -534 -1198
rect -526 -1206 -524 -1198
rect -510 -1206 -508 -1198
rect -356 -1206 -354 -1198
rect -346 -1206 -344 -1198
rect -330 -1206 -328 -1198
rect -145 -1206 -143 -1198
rect -135 -1206 -133 -1198
rect -119 -1206 -117 -1198
rect -860 -1424 -858 -1416
rect -852 -1424 -850 -1416
rect -846 -1424 -844 -1416
rect -838 -1424 -836 -1416
rect -830 -1424 -828 -1416
rect -822 -1424 -820 -1416
rect -816 -1424 -814 -1416
rect -810 -1424 -808 -1416
rect -799 -1424 -797 -1416
rect -786 -1424 -784 -1416
rect -778 -1424 -776 -1416
rect -770 -1424 -768 -1416
rect -758 -1424 -756 -1416
rect -739 -1424 -737 -1416
rect -634 -1424 -632 -1416
rect -626 -1424 -624 -1416
rect -620 -1424 -618 -1416
rect -612 -1424 -610 -1416
rect -604 -1424 -602 -1416
rect -596 -1424 -594 -1416
rect -590 -1424 -588 -1416
rect -584 -1424 -582 -1416
rect -573 -1424 -571 -1416
rect -560 -1424 -558 -1416
rect -552 -1424 -550 -1416
rect -544 -1424 -542 -1416
rect -532 -1424 -530 -1416
rect -513 -1424 -511 -1416
rect -416 -1424 -414 -1416
rect -408 -1424 -406 -1416
rect -402 -1424 -400 -1416
rect -394 -1424 -392 -1416
rect -386 -1424 -384 -1416
rect -378 -1424 -376 -1416
rect -372 -1424 -370 -1416
rect -366 -1424 -364 -1416
rect -355 -1424 -353 -1416
rect -342 -1424 -340 -1416
rect -334 -1424 -332 -1416
rect -326 -1424 -324 -1416
rect -314 -1424 -312 -1416
rect -295 -1424 -293 -1416
rect 18 -1417 20 -1409
rect 28 -1417 30 -1409
rect 44 -1417 46 -1409
rect -39 -1497 -37 -1489
rect 4 -1497 6 -1489
rect 14 -1497 16 -1489
rect 24 -1497 26 -1489
rect 33 -1497 35 -1489
rect -39 -1549 -37 -1541
<< ndiffusion >>
rect -304 -16 -303 -12
rect -301 -16 -300 -12
rect -330 -25 -329 -21
rect -327 -25 -319 -21
rect -317 -25 -316 -21
rect -183 -16 -182 -12
rect -180 -16 -179 -12
rect -209 -25 -208 -21
rect -206 -25 -198 -21
rect -196 -25 -195 -21
rect -69 -16 -68 -12
rect -66 -16 -65 -12
rect -95 -25 -94 -21
rect -92 -25 -84 -21
rect -82 -25 -81 -21
rect 31 -16 32 -12
rect 34 -16 35 -12
rect 5 -25 6 -21
rect 8 -25 16 -21
rect 18 -25 19 -21
rect -404 -234 -403 -230
rect -401 -234 -400 -230
rect -430 -243 -429 -239
rect -427 -243 -419 -239
rect -417 -243 -416 -239
rect -246 -234 -245 -230
rect -243 -234 -242 -230
rect -272 -243 -271 -239
rect -269 -243 -261 -239
rect -259 -243 -258 -239
rect -107 -234 -106 -230
rect -104 -234 -103 -230
rect -133 -243 -132 -239
rect -130 -243 -122 -239
rect -120 -243 -119 -239
rect 11 -234 12 -230
rect 14 -234 15 -230
rect -15 -243 -14 -239
rect -12 -243 -4 -239
rect -2 -243 -1 -239
rect -682 -402 -681 -398
rect -679 -402 -678 -398
rect -708 -411 -707 -407
rect -705 -411 -697 -407
rect -695 -411 -694 -407
rect -540 -432 -536 -420
rect -526 -432 -522 -420
rect -288 -432 -284 -420
rect -274 -432 -270 -420
rect 24 -402 25 -398
rect 27 -402 28 -398
rect -2 -411 -1 -407
rect 1 -411 9 -407
rect 11 -411 12 -407
rect -594 -436 -593 -432
rect -591 -436 -585 -432
rect -583 -436 -579 -432
rect -577 -436 -576 -432
rect -572 -436 -571 -432
rect -569 -436 -568 -432
rect -564 -436 -563 -432
rect -561 -436 -560 -432
rect -556 -436 -555 -432
rect -553 -436 -549 -432
rect -547 -436 -543 -432
rect -541 -436 -532 -432
rect -530 -436 -519 -432
rect -517 -436 -516 -432
rect -512 -436 -511 -432
rect -509 -436 -508 -432
rect -504 -436 -503 -432
rect -501 -436 -498 -432
rect -494 -436 -491 -432
rect -489 -436 -486 -432
rect -473 -436 -472 -432
rect -470 -436 -469 -432
rect -342 -436 -341 -432
rect -339 -436 -333 -432
rect -331 -436 -327 -432
rect -325 -436 -324 -432
rect -320 -436 -319 -432
rect -317 -436 -316 -432
rect -312 -436 -311 -432
rect -309 -436 -308 -432
rect -304 -436 -303 -432
rect -301 -436 -297 -432
rect -295 -436 -291 -432
rect -289 -436 -280 -432
rect -278 -436 -267 -432
rect -265 -436 -264 -432
rect -260 -436 -259 -432
rect -257 -436 -256 -432
rect -252 -436 -251 -432
rect -249 -436 -246 -432
rect -242 -436 -239 -432
rect -237 -436 -234 -432
rect -221 -436 -220 -432
rect -218 -436 -217 -432
rect -590 -443 -586 -436
rect -338 -443 -334 -436
rect -765 -481 -764 -477
rect -762 -481 -761 -477
rect -590 -449 -586 -445
rect -338 -449 -334 -445
rect -59 -481 -58 -477
rect -56 -481 -55 -477
rect -765 -533 -764 -529
rect -762 -533 -761 -529
rect -723 -533 -720 -529
rect -718 -533 -711 -529
rect -709 -533 -707 -529
rect -703 -533 -702 -529
rect -700 -533 -692 -529
rect -690 -533 -689 -529
rect -59 -533 -58 -529
rect -56 -533 -55 -529
rect -17 -533 -14 -529
rect -12 -533 -5 -529
rect -3 -533 -1 -529
rect 3 -533 4 -529
rect 6 -533 14 -529
rect 16 -533 17 -529
rect -689 -720 -688 -716
rect -686 -720 -685 -716
rect -715 -729 -714 -725
rect -712 -729 -704 -725
rect -702 -729 -701 -725
rect -511 -720 -510 -716
rect -508 -720 -507 -716
rect -537 -729 -536 -725
rect -534 -729 -526 -725
rect -524 -729 -523 -725
rect -331 -720 -330 -716
rect -328 -720 -327 -716
rect -357 -729 -356 -725
rect -354 -729 -346 -725
rect -344 -729 -343 -725
rect -120 -720 -119 -716
rect -117 -720 -116 -716
rect -146 -729 -145 -725
rect -143 -729 -135 -725
rect -133 -729 -132 -725
rect -762 -902 -758 -890
rect -748 -902 -744 -890
rect -536 -902 -532 -890
rect -522 -902 -518 -890
rect -318 -902 -314 -890
rect -304 -902 -300 -890
rect 43 -872 44 -868
rect 46 -872 47 -868
rect 17 -881 18 -877
rect 20 -881 28 -877
rect 30 -881 31 -877
rect -816 -906 -815 -902
rect -813 -906 -807 -902
rect -805 -906 -801 -902
rect -799 -906 -798 -902
rect -794 -906 -793 -902
rect -791 -906 -790 -902
rect -786 -906 -785 -902
rect -783 -906 -782 -902
rect -778 -906 -777 -902
rect -775 -906 -771 -902
rect -769 -906 -765 -902
rect -763 -906 -754 -902
rect -752 -906 -741 -902
rect -739 -906 -738 -902
rect -734 -906 -733 -902
rect -731 -906 -730 -902
rect -726 -906 -725 -902
rect -723 -906 -720 -902
rect -716 -906 -713 -902
rect -711 -906 -708 -902
rect -695 -906 -694 -902
rect -692 -906 -691 -902
rect -590 -906 -589 -902
rect -587 -906 -581 -902
rect -579 -906 -575 -902
rect -573 -906 -572 -902
rect -568 -906 -567 -902
rect -565 -906 -564 -902
rect -560 -906 -559 -902
rect -557 -906 -556 -902
rect -552 -906 -551 -902
rect -549 -906 -545 -902
rect -543 -906 -539 -902
rect -537 -906 -528 -902
rect -526 -906 -515 -902
rect -513 -906 -512 -902
rect -508 -906 -507 -902
rect -505 -906 -504 -902
rect -500 -906 -499 -902
rect -497 -906 -494 -902
rect -490 -906 -487 -902
rect -485 -906 -482 -902
rect -469 -906 -468 -902
rect -466 -906 -465 -902
rect -372 -906 -371 -902
rect -369 -906 -363 -902
rect -361 -906 -357 -902
rect -355 -906 -354 -902
rect -350 -906 -349 -902
rect -347 -906 -346 -902
rect -342 -906 -341 -902
rect -339 -906 -338 -902
rect -334 -906 -333 -902
rect -331 -906 -327 -902
rect -325 -906 -321 -902
rect -319 -906 -310 -902
rect -308 -906 -297 -902
rect -295 -906 -294 -902
rect -290 -906 -289 -902
rect -287 -906 -286 -902
rect -282 -906 -281 -902
rect -279 -906 -276 -902
rect -272 -906 -269 -902
rect -267 -906 -264 -902
rect -251 -906 -250 -902
rect -248 -906 -247 -902
rect -812 -913 -808 -906
rect -586 -913 -582 -906
rect -368 -913 -364 -906
rect -812 -919 -808 -915
rect -586 -919 -582 -915
rect -368 -919 -364 -915
rect -40 -951 -39 -947
rect -37 -951 -36 -947
rect -40 -1003 -39 -999
rect -37 -1003 -36 -999
rect 2 -1003 5 -999
rect 7 -1003 14 -999
rect 16 -1003 18 -999
rect 22 -1003 23 -999
rect 25 -1003 33 -999
rect 35 -1003 36 -999
rect -689 -1225 -688 -1221
rect -686 -1225 -685 -1221
rect -715 -1234 -714 -1230
rect -712 -1234 -704 -1230
rect -702 -1234 -701 -1230
rect -511 -1225 -510 -1221
rect -508 -1225 -507 -1221
rect -537 -1234 -536 -1230
rect -534 -1234 -526 -1230
rect -524 -1234 -523 -1230
rect -331 -1225 -330 -1221
rect -328 -1225 -327 -1221
rect -357 -1234 -356 -1230
rect -354 -1234 -346 -1230
rect -344 -1234 -343 -1230
rect -120 -1225 -119 -1221
rect -117 -1225 -116 -1221
rect -146 -1234 -145 -1230
rect -143 -1234 -135 -1230
rect -133 -1234 -132 -1230
rect -807 -1467 -803 -1455
rect -793 -1467 -789 -1455
rect -581 -1467 -577 -1455
rect -567 -1467 -563 -1455
rect -363 -1467 -359 -1455
rect -349 -1467 -345 -1455
rect 43 -1436 44 -1432
rect 46 -1436 47 -1432
rect 17 -1445 18 -1441
rect 20 -1445 28 -1441
rect 30 -1445 31 -1441
rect -861 -1471 -860 -1467
rect -858 -1471 -852 -1467
rect -850 -1471 -846 -1467
rect -844 -1471 -843 -1467
rect -839 -1471 -838 -1467
rect -836 -1471 -835 -1467
rect -831 -1471 -830 -1467
rect -828 -1471 -827 -1467
rect -823 -1471 -822 -1467
rect -820 -1471 -816 -1467
rect -814 -1471 -810 -1467
rect -808 -1471 -799 -1467
rect -797 -1471 -786 -1467
rect -784 -1471 -783 -1467
rect -779 -1471 -778 -1467
rect -776 -1471 -775 -1467
rect -771 -1471 -770 -1467
rect -768 -1471 -765 -1467
rect -761 -1471 -758 -1467
rect -756 -1471 -753 -1467
rect -740 -1471 -739 -1467
rect -737 -1471 -736 -1467
rect -635 -1471 -634 -1467
rect -632 -1471 -626 -1467
rect -624 -1471 -620 -1467
rect -618 -1471 -617 -1467
rect -613 -1471 -612 -1467
rect -610 -1471 -609 -1467
rect -605 -1471 -604 -1467
rect -602 -1471 -601 -1467
rect -597 -1471 -596 -1467
rect -594 -1471 -590 -1467
rect -588 -1471 -584 -1467
rect -582 -1471 -573 -1467
rect -571 -1471 -560 -1467
rect -558 -1471 -557 -1467
rect -553 -1471 -552 -1467
rect -550 -1471 -549 -1467
rect -545 -1471 -544 -1467
rect -542 -1471 -539 -1467
rect -535 -1471 -532 -1467
rect -530 -1471 -527 -1467
rect -514 -1471 -513 -1467
rect -511 -1471 -510 -1467
rect -417 -1471 -416 -1467
rect -414 -1471 -408 -1467
rect -406 -1471 -402 -1467
rect -400 -1471 -399 -1467
rect -395 -1471 -394 -1467
rect -392 -1471 -391 -1467
rect -387 -1471 -386 -1467
rect -384 -1471 -383 -1467
rect -379 -1471 -378 -1467
rect -376 -1471 -372 -1467
rect -370 -1471 -366 -1467
rect -364 -1471 -355 -1467
rect -353 -1471 -342 -1467
rect -340 -1471 -339 -1467
rect -335 -1471 -334 -1467
rect -332 -1471 -331 -1467
rect -327 -1471 -326 -1467
rect -324 -1471 -321 -1467
rect -317 -1471 -314 -1467
rect -312 -1471 -309 -1467
rect -296 -1471 -295 -1467
rect -293 -1471 -292 -1467
rect -857 -1478 -853 -1471
rect -631 -1478 -627 -1471
rect -413 -1478 -409 -1471
rect -857 -1484 -853 -1480
rect -631 -1484 -627 -1480
rect -413 -1484 -409 -1480
rect -40 -1515 -39 -1511
rect -37 -1515 -36 -1511
rect -40 -1567 -39 -1563
rect -37 -1567 -36 -1563
rect 2 -1567 5 -1563
rect 7 -1567 14 -1563
rect 16 -1567 18 -1563
rect 22 -1567 23 -1563
rect 25 -1567 33 -1563
rect 35 -1567 36 -1563
<< pdiffusion >>
rect -330 3 -329 11
rect -327 3 -324 11
rect -320 3 -319 11
rect -317 3 -316 11
rect -304 3 -303 11
rect -301 3 -300 11
rect -209 3 -208 11
rect -206 3 -203 11
rect -199 3 -198 11
rect -196 3 -195 11
rect -183 3 -182 11
rect -180 3 -179 11
rect -95 3 -94 11
rect -92 3 -89 11
rect -85 3 -84 11
rect -82 3 -81 11
rect -69 3 -68 11
rect -66 3 -65 11
rect 5 3 6 11
rect 8 3 11 11
rect 15 3 16 11
rect 18 3 19 11
rect 31 3 32 11
rect 34 3 35 11
rect -430 -215 -429 -207
rect -427 -215 -424 -207
rect -420 -215 -419 -207
rect -417 -215 -416 -207
rect -404 -215 -403 -207
rect -401 -215 -400 -207
rect -272 -215 -271 -207
rect -269 -215 -266 -207
rect -262 -215 -261 -207
rect -259 -215 -258 -207
rect -246 -215 -245 -207
rect -243 -215 -242 -207
rect -133 -215 -132 -207
rect -130 -215 -127 -207
rect -123 -215 -122 -207
rect -120 -215 -119 -207
rect -107 -215 -106 -207
rect -104 -215 -103 -207
rect -15 -215 -14 -207
rect -12 -215 -9 -207
rect -5 -215 -4 -207
rect -2 -215 -1 -207
rect 11 -215 12 -207
rect 14 -215 15 -207
rect -708 -383 -707 -375
rect -705 -383 -702 -375
rect -698 -383 -697 -375
rect -695 -383 -694 -375
rect -682 -383 -681 -375
rect -679 -383 -678 -375
rect -590 -381 -586 -370
rect -338 -381 -334 -370
rect -594 -389 -593 -381
rect -591 -389 -585 -381
rect -583 -389 -579 -381
rect -577 -389 -576 -381
rect -572 -389 -571 -381
rect -569 -389 -568 -381
rect -564 -389 -563 -381
rect -561 -389 -560 -381
rect -556 -389 -555 -381
rect -553 -389 -549 -381
rect -547 -389 -543 -381
rect -541 -389 -540 -381
rect -536 -389 -532 -381
rect -530 -389 -526 -381
rect -522 -389 -519 -381
rect -517 -389 -516 -381
rect -512 -389 -511 -381
rect -509 -389 -508 -381
rect -504 -389 -503 -381
rect -501 -389 -498 -381
rect -494 -389 -491 -381
rect -489 -389 -486 -381
rect -473 -389 -472 -381
rect -470 -389 -469 -381
rect -342 -389 -341 -381
rect -339 -389 -333 -381
rect -331 -389 -327 -381
rect -325 -389 -324 -381
rect -320 -389 -319 -381
rect -317 -389 -316 -381
rect -312 -389 -311 -381
rect -309 -389 -308 -381
rect -304 -389 -303 -381
rect -301 -389 -297 -381
rect -295 -389 -291 -381
rect -289 -389 -288 -381
rect -284 -389 -280 -381
rect -278 -389 -274 -381
rect -270 -389 -267 -381
rect -265 -389 -264 -381
rect -260 -389 -259 -381
rect -257 -389 -256 -381
rect -252 -389 -251 -381
rect -249 -389 -246 -381
rect -242 -389 -239 -381
rect -237 -389 -234 -381
rect -221 -389 -220 -381
rect -218 -389 -217 -381
rect -2 -383 -1 -375
rect 1 -383 4 -375
rect 8 -383 9 -375
rect 11 -383 12 -375
rect 24 -383 25 -375
rect 27 -383 28 -375
rect -765 -463 -764 -455
rect -762 -463 -761 -455
rect -723 -463 -721 -455
rect -719 -463 -711 -455
rect -709 -463 -707 -455
rect -703 -463 -701 -455
rect -699 -463 -692 -455
rect -690 -463 -689 -455
rect -765 -515 -764 -507
rect -762 -515 -761 -507
rect -59 -463 -58 -455
rect -56 -463 -55 -455
rect -17 -463 -15 -455
rect -13 -463 -5 -455
rect -3 -463 -1 -455
rect 3 -463 5 -455
rect 7 -463 14 -455
rect 16 -463 17 -455
rect -59 -515 -58 -507
rect -56 -515 -55 -507
rect -715 -701 -714 -693
rect -712 -701 -709 -693
rect -705 -701 -704 -693
rect -702 -701 -701 -693
rect -689 -701 -688 -693
rect -686 -701 -685 -693
rect -537 -701 -536 -693
rect -534 -701 -531 -693
rect -527 -701 -526 -693
rect -524 -701 -523 -693
rect -511 -701 -510 -693
rect -508 -701 -507 -693
rect -357 -701 -356 -693
rect -354 -701 -351 -693
rect -347 -701 -346 -693
rect -344 -701 -343 -693
rect -331 -701 -330 -693
rect -328 -701 -327 -693
rect -146 -701 -145 -693
rect -143 -701 -140 -693
rect -136 -701 -135 -693
rect -133 -701 -132 -693
rect -120 -701 -119 -693
rect -117 -701 -116 -693
rect -812 -851 -808 -840
rect -586 -851 -582 -840
rect -368 -851 -364 -840
rect -816 -859 -815 -851
rect -813 -859 -807 -851
rect -805 -859 -801 -851
rect -799 -859 -798 -851
rect -794 -859 -793 -851
rect -791 -859 -790 -851
rect -786 -859 -785 -851
rect -783 -859 -782 -851
rect -778 -859 -777 -851
rect -775 -859 -771 -851
rect -769 -859 -765 -851
rect -763 -859 -762 -851
rect -758 -859 -754 -851
rect -752 -859 -748 -851
rect -744 -859 -741 -851
rect -739 -859 -738 -851
rect -734 -859 -733 -851
rect -731 -859 -730 -851
rect -726 -859 -725 -851
rect -723 -859 -720 -851
rect -716 -859 -713 -851
rect -711 -859 -708 -851
rect -695 -859 -694 -851
rect -692 -859 -691 -851
rect -590 -859 -589 -851
rect -587 -859 -581 -851
rect -579 -859 -575 -851
rect -573 -859 -572 -851
rect -568 -859 -567 -851
rect -565 -859 -564 -851
rect -560 -859 -559 -851
rect -557 -859 -556 -851
rect -552 -859 -551 -851
rect -549 -859 -545 -851
rect -543 -859 -539 -851
rect -537 -859 -536 -851
rect -532 -859 -528 -851
rect -526 -859 -522 -851
rect -518 -859 -515 -851
rect -513 -859 -512 -851
rect -508 -859 -507 -851
rect -505 -859 -504 -851
rect -500 -859 -499 -851
rect -497 -859 -494 -851
rect -490 -859 -487 -851
rect -485 -859 -482 -851
rect -469 -859 -468 -851
rect -466 -859 -465 -851
rect -372 -859 -371 -851
rect -369 -859 -363 -851
rect -361 -859 -357 -851
rect -355 -859 -354 -851
rect -350 -859 -349 -851
rect -347 -859 -346 -851
rect -342 -859 -341 -851
rect -339 -859 -338 -851
rect -334 -859 -333 -851
rect -331 -859 -327 -851
rect -325 -859 -321 -851
rect -319 -859 -318 -851
rect -314 -859 -310 -851
rect -308 -859 -304 -851
rect -300 -859 -297 -851
rect -295 -859 -294 -851
rect -290 -859 -289 -851
rect -287 -859 -286 -851
rect -282 -859 -281 -851
rect -279 -859 -276 -851
rect -272 -859 -269 -851
rect -267 -859 -264 -851
rect -251 -859 -250 -851
rect -248 -859 -247 -851
rect 17 -853 18 -845
rect 20 -853 23 -845
rect 27 -853 28 -845
rect 30 -853 31 -845
rect 43 -853 44 -845
rect 46 -853 47 -845
rect -40 -933 -39 -925
rect -37 -933 -36 -925
rect 2 -933 4 -925
rect 6 -933 14 -925
rect 16 -933 18 -925
rect 22 -933 24 -925
rect 26 -933 33 -925
rect 35 -933 36 -925
rect -40 -985 -39 -977
rect -37 -985 -36 -977
rect -715 -1206 -714 -1198
rect -712 -1206 -709 -1198
rect -705 -1206 -704 -1198
rect -702 -1206 -701 -1198
rect -689 -1206 -688 -1198
rect -686 -1206 -685 -1198
rect -537 -1206 -536 -1198
rect -534 -1206 -531 -1198
rect -527 -1206 -526 -1198
rect -524 -1206 -523 -1198
rect -511 -1206 -510 -1198
rect -508 -1206 -507 -1198
rect -357 -1206 -356 -1198
rect -354 -1206 -351 -1198
rect -347 -1206 -346 -1198
rect -344 -1206 -343 -1198
rect -331 -1206 -330 -1198
rect -328 -1206 -327 -1198
rect -146 -1206 -145 -1198
rect -143 -1206 -140 -1198
rect -136 -1206 -135 -1198
rect -133 -1206 -132 -1198
rect -120 -1206 -119 -1198
rect -117 -1206 -116 -1198
rect -857 -1416 -853 -1405
rect -631 -1416 -627 -1405
rect -413 -1416 -409 -1405
rect -861 -1424 -860 -1416
rect -858 -1424 -852 -1416
rect -850 -1424 -846 -1416
rect -844 -1424 -843 -1416
rect -839 -1424 -838 -1416
rect -836 -1424 -835 -1416
rect -831 -1424 -830 -1416
rect -828 -1424 -827 -1416
rect -823 -1424 -822 -1416
rect -820 -1424 -816 -1416
rect -814 -1424 -810 -1416
rect -808 -1424 -807 -1416
rect -803 -1424 -799 -1416
rect -797 -1424 -793 -1416
rect -789 -1424 -786 -1416
rect -784 -1424 -783 -1416
rect -779 -1424 -778 -1416
rect -776 -1424 -775 -1416
rect -771 -1424 -770 -1416
rect -768 -1424 -765 -1416
rect -761 -1424 -758 -1416
rect -756 -1424 -753 -1416
rect -740 -1424 -739 -1416
rect -737 -1424 -736 -1416
rect -635 -1424 -634 -1416
rect -632 -1424 -626 -1416
rect -624 -1424 -620 -1416
rect -618 -1424 -617 -1416
rect -613 -1424 -612 -1416
rect -610 -1424 -609 -1416
rect -605 -1424 -604 -1416
rect -602 -1424 -601 -1416
rect -597 -1424 -596 -1416
rect -594 -1424 -590 -1416
rect -588 -1424 -584 -1416
rect -582 -1424 -581 -1416
rect -577 -1424 -573 -1416
rect -571 -1424 -567 -1416
rect -563 -1424 -560 -1416
rect -558 -1424 -557 -1416
rect -553 -1424 -552 -1416
rect -550 -1424 -549 -1416
rect -545 -1424 -544 -1416
rect -542 -1424 -539 -1416
rect -535 -1424 -532 -1416
rect -530 -1424 -527 -1416
rect -514 -1424 -513 -1416
rect -511 -1424 -510 -1416
rect -417 -1424 -416 -1416
rect -414 -1424 -408 -1416
rect -406 -1424 -402 -1416
rect -400 -1424 -399 -1416
rect -395 -1424 -394 -1416
rect -392 -1424 -391 -1416
rect -387 -1424 -386 -1416
rect -384 -1424 -383 -1416
rect -379 -1424 -378 -1416
rect -376 -1424 -372 -1416
rect -370 -1424 -366 -1416
rect -364 -1424 -363 -1416
rect -359 -1424 -355 -1416
rect -353 -1424 -349 -1416
rect -345 -1424 -342 -1416
rect -340 -1424 -339 -1416
rect -335 -1424 -334 -1416
rect -332 -1424 -331 -1416
rect -327 -1424 -326 -1416
rect -324 -1424 -321 -1416
rect -317 -1424 -314 -1416
rect -312 -1424 -309 -1416
rect -296 -1424 -295 -1416
rect -293 -1424 -292 -1416
rect 17 -1417 18 -1409
rect 20 -1417 23 -1409
rect 27 -1417 28 -1409
rect 30 -1417 31 -1409
rect 43 -1417 44 -1409
rect 46 -1417 47 -1409
rect -40 -1497 -39 -1489
rect -37 -1497 -36 -1489
rect 2 -1497 4 -1489
rect 6 -1497 14 -1489
rect 16 -1497 18 -1489
rect 22 -1497 24 -1489
rect 26 -1497 33 -1489
rect 35 -1497 36 -1489
rect -40 -1549 -39 -1541
rect -37 -1549 -36 -1541
<< ndcontact >>
rect -308 -16 -304 -12
rect -300 -16 -296 -12
rect -334 -25 -330 -21
rect -316 -25 -312 -21
rect -187 -16 -183 -12
rect -179 -16 -175 -12
rect -213 -25 -209 -21
rect -195 -25 -191 -21
rect -73 -16 -69 -12
rect -65 -16 -61 -12
rect -99 -25 -95 -21
rect -81 -25 -77 -21
rect 27 -16 31 -12
rect 35 -16 39 -12
rect 1 -25 5 -21
rect 19 -25 23 -21
rect -408 -234 -404 -230
rect -400 -234 -396 -230
rect -434 -243 -430 -239
rect -416 -243 -412 -239
rect -250 -234 -246 -230
rect -242 -234 -238 -230
rect -276 -243 -272 -239
rect -258 -243 -254 -239
rect -111 -234 -107 -230
rect -103 -234 -99 -230
rect -137 -243 -133 -239
rect -119 -243 -115 -239
rect 7 -234 11 -230
rect 15 -234 19 -230
rect -19 -243 -15 -239
rect -1 -243 3 -239
rect -686 -402 -682 -398
rect -678 -402 -674 -398
rect -712 -411 -708 -407
rect -694 -411 -690 -407
rect -540 -420 -536 -416
rect -526 -420 -522 -416
rect -288 -420 -284 -416
rect -274 -420 -270 -416
rect 20 -402 24 -398
rect 28 -402 32 -398
rect -6 -411 -2 -407
rect 12 -411 16 -407
rect -598 -436 -594 -432
rect -576 -436 -572 -432
rect -568 -436 -564 -432
rect -560 -436 -556 -432
rect -516 -436 -512 -432
rect -508 -436 -504 -432
rect -498 -436 -494 -432
rect -486 -436 -482 -432
rect -477 -436 -473 -432
rect -469 -436 -465 -432
rect -346 -436 -342 -432
rect -324 -436 -320 -432
rect -316 -436 -312 -432
rect -308 -436 -304 -432
rect -264 -436 -260 -432
rect -256 -436 -252 -432
rect -246 -436 -242 -432
rect -234 -436 -230 -432
rect -225 -436 -221 -432
rect -217 -436 -213 -432
rect -769 -481 -765 -477
rect -761 -481 -757 -477
rect -590 -453 -586 -449
rect -338 -453 -334 -449
rect -63 -481 -59 -477
rect -55 -481 -51 -477
rect -769 -533 -765 -529
rect -761 -533 -757 -529
rect -727 -533 -723 -529
rect -707 -533 -703 -529
rect -689 -533 -685 -529
rect -63 -533 -59 -529
rect -55 -533 -51 -529
rect -21 -533 -17 -529
rect -1 -533 3 -529
rect 17 -533 21 -529
rect -693 -720 -689 -716
rect -685 -720 -681 -716
rect -719 -729 -715 -725
rect -701 -729 -697 -725
rect -515 -720 -511 -716
rect -507 -720 -503 -716
rect -541 -729 -537 -725
rect -523 -729 -519 -725
rect -335 -720 -331 -716
rect -327 -720 -323 -716
rect -361 -729 -357 -725
rect -343 -729 -339 -725
rect -124 -720 -120 -716
rect -116 -720 -112 -716
rect -150 -729 -146 -725
rect -132 -729 -128 -725
rect -762 -890 -758 -886
rect -748 -890 -744 -886
rect -536 -890 -532 -886
rect -522 -890 -518 -886
rect -318 -890 -314 -886
rect -304 -890 -300 -886
rect 39 -872 43 -868
rect 47 -872 51 -868
rect 13 -881 17 -877
rect 31 -881 35 -877
rect -820 -906 -816 -902
rect -798 -906 -794 -902
rect -790 -906 -786 -902
rect -782 -906 -778 -902
rect -738 -906 -734 -902
rect -730 -906 -726 -902
rect -720 -906 -716 -902
rect -708 -906 -704 -902
rect -699 -906 -695 -902
rect -691 -906 -687 -902
rect -594 -906 -590 -902
rect -572 -906 -568 -902
rect -564 -906 -560 -902
rect -556 -906 -552 -902
rect -512 -906 -508 -902
rect -504 -906 -500 -902
rect -494 -906 -490 -902
rect -482 -906 -478 -902
rect -473 -906 -469 -902
rect -465 -906 -461 -902
rect -376 -906 -372 -902
rect -354 -906 -350 -902
rect -346 -906 -342 -902
rect -338 -906 -334 -902
rect -294 -906 -290 -902
rect -286 -906 -282 -902
rect -276 -906 -272 -902
rect -264 -906 -260 -902
rect -255 -906 -251 -902
rect -247 -906 -243 -902
rect -812 -923 -808 -919
rect -586 -923 -582 -919
rect -368 -923 -364 -919
rect -44 -951 -40 -947
rect -36 -951 -32 -947
rect -44 -1003 -40 -999
rect -36 -1003 -32 -999
rect -2 -1003 2 -999
rect 18 -1003 22 -999
rect 36 -1003 40 -999
rect -693 -1225 -689 -1221
rect -685 -1225 -681 -1221
rect -719 -1234 -715 -1230
rect -701 -1234 -697 -1230
rect -515 -1225 -511 -1221
rect -507 -1225 -503 -1221
rect -541 -1234 -537 -1230
rect -523 -1234 -519 -1230
rect -335 -1225 -331 -1221
rect -327 -1225 -323 -1221
rect -361 -1234 -357 -1230
rect -343 -1234 -339 -1230
rect -124 -1225 -120 -1221
rect -116 -1225 -112 -1221
rect -150 -1234 -146 -1230
rect -132 -1234 -128 -1230
rect -807 -1455 -803 -1451
rect -793 -1455 -789 -1451
rect -581 -1455 -577 -1451
rect -567 -1455 -563 -1451
rect -363 -1455 -359 -1451
rect -349 -1455 -345 -1451
rect 39 -1436 43 -1432
rect 47 -1436 51 -1432
rect 13 -1445 17 -1441
rect 31 -1445 35 -1441
rect -865 -1471 -861 -1467
rect -843 -1471 -839 -1467
rect -835 -1471 -831 -1467
rect -827 -1471 -823 -1467
rect -783 -1471 -779 -1467
rect -775 -1471 -771 -1467
rect -765 -1471 -761 -1467
rect -753 -1471 -749 -1467
rect -744 -1471 -740 -1467
rect -736 -1471 -732 -1467
rect -639 -1471 -635 -1467
rect -617 -1471 -613 -1467
rect -609 -1471 -605 -1467
rect -601 -1471 -597 -1467
rect -557 -1471 -553 -1467
rect -549 -1471 -545 -1467
rect -539 -1471 -535 -1467
rect -527 -1471 -523 -1467
rect -518 -1471 -514 -1467
rect -510 -1471 -506 -1467
rect -421 -1471 -417 -1467
rect -399 -1471 -395 -1467
rect -391 -1471 -387 -1467
rect -383 -1471 -379 -1467
rect -339 -1471 -335 -1467
rect -331 -1471 -327 -1467
rect -321 -1471 -317 -1467
rect -309 -1471 -305 -1467
rect -300 -1471 -296 -1467
rect -292 -1471 -288 -1467
rect -857 -1488 -853 -1484
rect -631 -1488 -627 -1484
rect -413 -1488 -409 -1484
rect -44 -1515 -40 -1511
rect -36 -1515 -32 -1511
rect -44 -1567 -40 -1563
rect -36 -1567 -32 -1563
rect -2 -1567 2 -1563
rect 18 -1567 22 -1563
rect 36 -1567 40 -1563
<< pdcontact >>
rect -334 3 -330 11
rect -324 3 -320 11
rect -316 3 -312 11
rect -308 3 -304 11
rect -300 3 -296 11
rect -213 3 -209 11
rect -203 3 -199 11
rect -195 3 -191 11
rect -187 3 -183 11
rect -179 3 -175 11
rect -99 3 -95 11
rect -89 3 -85 11
rect -81 3 -77 11
rect -73 3 -69 11
rect -65 3 -61 11
rect 1 3 5 11
rect 11 3 15 11
rect 19 3 23 11
rect 27 3 31 11
rect 35 3 39 11
rect -434 -215 -430 -207
rect -424 -215 -420 -207
rect -416 -215 -412 -207
rect -408 -215 -404 -207
rect -400 -215 -396 -207
rect -276 -215 -272 -207
rect -266 -215 -262 -207
rect -258 -215 -254 -207
rect -250 -215 -246 -207
rect -242 -215 -238 -207
rect -137 -215 -133 -207
rect -127 -215 -123 -207
rect -119 -215 -115 -207
rect -111 -215 -107 -207
rect -103 -215 -99 -207
rect -19 -215 -15 -207
rect -9 -215 -5 -207
rect -1 -215 3 -207
rect 7 -215 11 -207
rect 15 -215 19 -207
rect -590 -370 -586 -366
rect -712 -383 -708 -375
rect -702 -383 -698 -375
rect -694 -383 -690 -375
rect -686 -383 -682 -375
rect -678 -383 -674 -375
rect -338 -370 -334 -366
rect -598 -389 -594 -381
rect -576 -389 -572 -381
rect -568 -389 -564 -381
rect -560 -389 -556 -381
rect -540 -389 -536 -381
rect -526 -389 -522 -381
rect -516 -389 -512 -381
rect -508 -389 -504 -381
rect -498 -389 -494 -381
rect -486 -389 -482 -381
rect -477 -389 -473 -381
rect -469 -389 -465 -381
rect -346 -389 -342 -381
rect -324 -389 -320 -381
rect -316 -389 -312 -381
rect -308 -389 -304 -381
rect -288 -389 -284 -381
rect -274 -389 -270 -381
rect -264 -389 -260 -381
rect -256 -389 -252 -381
rect -246 -389 -242 -381
rect -234 -389 -230 -381
rect -225 -389 -221 -381
rect -217 -389 -213 -381
rect -6 -383 -2 -375
rect 4 -383 8 -375
rect 12 -383 16 -375
rect 20 -383 24 -375
rect 28 -383 32 -375
rect -769 -463 -765 -455
rect -761 -463 -757 -455
rect -727 -463 -723 -455
rect -707 -463 -703 -455
rect -689 -463 -685 -455
rect -769 -515 -765 -507
rect -761 -515 -757 -507
rect -63 -463 -59 -455
rect -55 -463 -51 -455
rect -21 -463 -17 -455
rect -1 -463 3 -455
rect 17 -463 21 -455
rect -63 -515 -59 -507
rect -55 -515 -51 -507
rect -719 -701 -715 -693
rect -709 -701 -705 -693
rect -701 -701 -697 -693
rect -693 -701 -689 -693
rect -685 -701 -681 -693
rect -541 -701 -537 -693
rect -531 -701 -527 -693
rect -523 -701 -519 -693
rect -515 -701 -511 -693
rect -507 -701 -503 -693
rect -361 -701 -357 -693
rect -351 -701 -347 -693
rect -343 -701 -339 -693
rect -335 -701 -331 -693
rect -327 -701 -323 -693
rect -150 -701 -146 -693
rect -140 -701 -136 -693
rect -132 -701 -128 -693
rect -124 -701 -120 -693
rect -116 -701 -112 -693
rect -812 -840 -808 -836
rect -586 -840 -582 -836
rect -368 -840 -364 -836
rect -820 -859 -816 -851
rect -798 -859 -794 -851
rect -790 -859 -786 -851
rect -782 -859 -778 -851
rect -762 -859 -758 -851
rect -748 -859 -744 -851
rect -738 -859 -734 -851
rect -730 -859 -726 -851
rect -720 -859 -716 -851
rect -708 -859 -704 -851
rect -699 -859 -695 -851
rect -691 -859 -687 -851
rect -594 -859 -590 -851
rect -572 -859 -568 -851
rect -564 -859 -560 -851
rect -556 -859 -552 -851
rect -536 -859 -532 -851
rect -522 -859 -518 -851
rect -512 -859 -508 -851
rect -504 -859 -500 -851
rect -494 -859 -490 -851
rect -482 -859 -478 -851
rect -473 -859 -469 -851
rect -465 -859 -461 -851
rect -376 -859 -372 -851
rect -354 -859 -350 -851
rect -346 -859 -342 -851
rect -338 -859 -334 -851
rect -318 -859 -314 -851
rect -304 -859 -300 -851
rect -294 -859 -290 -851
rect -286 -859 -282 -851
rect -276 -859 -272 -851
rect -264 -859 -260 -851
rect -255 -859 -251 -851
rect -247 -859 -243 -851
rect 13 -853 17 -845
rect 23 -853 27 -845
rect 31 -853 35 -845
rect 39 -853 43 -845
rect 47 -853 51 -845
rect -44 -933 -40 -925
rect -36 -933 -32 -925
rect -2 -933 2 -925
rect 18 -933 22 -925
rect 36 -933 40 -925
rect -44 -985 -40 -977
rect -36 -985 -32 -977
rect -719 -1206 -715 -1198
rect -709 -1206 -705 -1198
rect -701 -1206 -697 -1198
rect -693 -1206 -689 -1198
rect -685 -1206 -681 -1198
rect -541 -1206 -537 -1198
rect -531 -1206 -527 -1198
rect -523 -1206 -519 -1198
rect -515 -1206 -511 -1198
rect -507 -1206 -503 -1198
rect -361 -1206 -357 -1198
rect -351 -1206 -347 -1198
rect -343 -1206 -339 -1198
rect -335 -1206 -331 -1198
rect -327 -1206 -323 -1198
rect -150 -1206 -146 -1198
rect -140 -1206 -136 -1198
rect -132 -1206 -128 -1198
rect -124 -1206 -120 -1198
rect -116 -1206 -112 -1198
rect -857 -1405 -853 -1401
rect -631 -1405 -627 -1401
rect -413 -1405 -409 -1401
rect -865 -1424 -861 -1416
rect -843 -1424 -839 -1416
rect -835 -1424 -831 -1416
rect -827 -1424 -823 -1416
rect -807 -1424 -803 -1416
rect -793 -1424 -789 -1416
rect -783 -1424 -779 -1416
rect -775 -1424 -771 -1416
rect -765 -1424 -761 -1416
rect -753 -1424 -749 -1416
rect -744 -1424 -740 -1416
rect -736 -1424 -732 -1416
rect -639 -1424 -635 -1416
rect -617 -1424 -613 -1416
rect -609 -1424 -605 -1416
rect -601 -1424 -597 -1416
rect -581 -1424 -577 -1416
rect -567 -1424 -563 -1416
rect -557 -1424 -553 -1416
rect -549 -1424 -545 -1416
rect -539 -1424 -535 -1416
rect -527 -1424 -523 -1416
rect -518 -1424 -514 -1416
rect -510 -1424 -506 -1416
rect -421 -1424 -417 -1416
rect -399 -1424 -395 -1416
rect -391 -1424 -387 -1416
rect -383 -1424 -379 -1416
rect -363 -1424 -359 -1416
rect -349 -1424 -345 -1416
rect -339 -1424 -335 -1416
rect -331 -1424 -327 -1416
rect -321 -1424 -317 -1416
rect -309 -1424 -305 -1416
rect -300 -1424 -296 -1416
rect -292 -1424 -288 -1416
rect 13 -1417 17 -1409
rect 23 -1417 27 -1409
rect 31 -1417 35 -1409
rect 39 -1417 43 -1409
rect 47 -1417 51 -1409
rect -44 -1497 -40 -1489
rect -36 -1497 -32 -1489
rect -2 -1497 2 -1489
rect 18 -1497 22 -1489
rect 36 -1497 40 -1489
rect -44 -1549 -40 -1541
rect -36 -1549 -32 -1541
<< polysilicon >>
rect -329 11 -327 14
rect -319 11 -317 14
rect -303 11 -301 14
rect -208 11 -206 14
rect -198 11 -196 14
rect -182 11 -180 14
rect -94 11 -92 14
rect -84 11 -82 14
rect -68 11 -66 14
rect 6 11 8 14
rect 16 11 18 14
rect 32 11 34 14
rect -329 -21 -327 3
rect -319 -21 -317 3
rect -303 -12 -301 3
rect -329 -28 -327 -25
rect -319 -28 -317 -25
rect -303 -28 -301 -16
rect -208 -21 -206 3
rect -198 -21 -196 3
rect -182 -12 -180 3
rect -208 -28 -206 -25
rect -198 -28 -196 -25
rect -182 -28 -180 -16
rect -94 -21 -92 3
rect -84 -21 -82 3
rect -68 -12 -66 3
rect -94 -28 -92 -25
rect -84 -28 -82 -25
rect -68 -28 -66 -16
rect 6 -21 8 3
rect 16 -21 18 3
rect 32 -12 34 3
rect 6 -28 8 -25
rect 16 -28 18 -25
rect 32 -28 34 -16
rect -429 -207 -427 -204
rect -419 -207 -417 -204
rect -403 -207 -401 -204
rect -271 -207 -269 -204
rect -261 -207 -259 -204
rect -245 -207 -243 -204
rect -132 -207 -130 -204
rect -122 -207 -120 -204
rect -106 -207 -104 -204
rect -14 -207 -12 -204
rect -4 -207 -2 -204
rect 12 -207 14 -204
rect -429 -239 -427 -215
rect -419 -239 -417 -215
rect -403 -230 -401 -215
rect -429 -246 -427 -243
rect -419 -246 -417 -243
rect -403 -246 -401 -234
rect -271 -239 -269 -215
rect -261 -239 -259 -215
rect -245 -230 -243 -215
rect -271 -246 -269 -243
rect -261 -246 -259 -243
rect -245 -246 -243 -234
rect -132 -239 -130 -215
rect -122 -239 -120 -215
rect -106 -230 -104 -215
rect -132 -246 -130 -243
rect -122 -246 -120 -243
rect -106 -246 -104 -234
rect -14 -239 -12 -215
rect -4 -239 -2 -215
rect 12 -230 14 -215
rect -14 -246 -12 -243
rect -4 -246 -2 -243
rect 12 -246 14 -234
rect -563 -368 -561 -358
rect -707 -375 -705 -372
rect -697 -375 -695 -372
rect -681 -375 -679 -372
rect -593 -381 -591 -378
rect -585 -370 -509 -368
rect -585 -381 -583 -370
rect -579 -375 -561 -373
rect -579 -381 -577 -375
rect -571 -381 -569 -378
rect -563 -381 -561 -375
rect -555 -381 -553 -378
rect -549 -381 -547 -370
rect -543 -381 -541 -378
rect -532 -381 -530 -378
rect -519 -381 -517 -378
rect -511 -381 -509 -370
rect -311 -368 -309 -358
rect -503 -381 -501 -378
rect -491 -381 -489 -377
rect -472 -381 -470 -378
rect -341 -381 -339 -378
rect -333 -370 -257 -368
rect -333 -381 -331 -370
rect -327 -375 -309 -373
rect -327 -381 -325 -375
rect -319 -381 -317 -378
rect -311 -381 -309 -375
rect -303 -381 -301 -378
rect -297 -381 -295 -370
rect -291 -381 -289 -378
rect -280 -381 -278 -378
rect -267 -381 -265 -378
rect -259 -381 -257 -370
rect -1 -375 1 -372
rect 9 -375 11 -372
rect 25 -375 27 -372
rect -251 -381 -249 -378
rect -239 -381 -237 -377
rect -220 -381 -218 -378
rect -707 -407 -705 -383
rect -697 -407 -695 -383
rect -681 -398 -679 -383
rect -593 -391 -591 -389
rect -585 -391 -583 -389
rect -593 -393 -583 -391
rect -707 -414 -705 -411
rect -697 -414 -695 -411
rect -681 -414 -679 -402
rect -593 -432 -591 -393
rect -585 -432 -583 -393
rect -579 -432 -577 -389
rect -571 -432 -569 -389
rect -563 -391 -561 -389
rect -555 -391 -553 -389
rect -563 -393 -553 -391
rect -563 -415 -561 -393
rect -563 -432 -561 -420
rect -555 -432 -553 -393
rect -549 -432 -547 -389
rect -543 -432 -541 -389
rect -532 -424 -530 -389
rect -532 -432 -530 -429
rect -519 -432 -517 -389
rect -511 -432 -509 -389
rect -503 -432 -501 -389
rect -491 -432 -489 -389
rect -472 -432 -470 -389
rect -341 -391 -339 -389
rect -333 -391 -331 -389
rect -341 -393 -331 -391
rect -341 -432 -339 -393
rect -333 -432 -331 -393
rect -327 -432 -325 -389
rect -319 -432 -317 -389
rect -311 -391 -309 -389
rect -303 -391 -301 -389
rect -311 -393 -301 -391
rect -311 -415 -309 -393
rect -311 -432 -309 -420
rect -303 -432 -301 -393
rect -297 -432 -295 -389
rect -291 -432 -289 -389
rect -280 -424 -278 -389
rect -280 -432 -278 -429
rect -267 -432 -265 -389
rect -259 -432 -257 -389
rect -251 -432 -249 -389
rect -239 -432 -237 -389
rect -220 -432 -218 -389
rect -1 -407 1 -383
rect 9 -407 11 -383
rect 25 -398 27 -383
rect -1 -414 1 -411
rect 9 -414 11 -411
rect 25 -414 27 -402
rect -602 -443 -600 -437
rect -593 -439 -591 -436
rect -585 -439 -583 -436
rect -579 -439 -577 -436
rect -571 -443 -569 -436
rect -563 -439 -561 -436
rect -555 -439 -553 -436
rect -549 -439 -547 -436
rect -543 -443 -541 -436
rect -532 -439 -530 -436
rect -519 -443 -517 -436
rect -511 -439 -509 -436
rect -503 -439 -501 -436
rect -491 -439 -489 -436
rect -472 -439 -470 -436
rect -721 -445 -681 -443
rect -602 -445 -590 -443
rect -586 -445 -517 -443
rect -350 -443 -348 -438
rect -341 -439 -339 -436
rect -333 -439 -331 -436
rect -327 -439 -325 -436
rect -319 -443 -317 -436
rect -311 -439 -309 -436
rect -303 -439 -301 -436
rect -297 -439 -295 -436
rect -291 -443 -289 -436
rect -280 -439 -278 -436
rect -267 -443 -265 -436
rect -259 -439 -257 -436
rect -251 -439 -249 -436
rect -239 -439 -237 -436
rect -220 -439 -218 -436
rect -350 -445 -338 -443
rect -334 -445 -265 -443
rect -15 -445 25 -443
rect -764 -455 -762 -452
rect -721 -455 -719 -445
rect -711 -455 -709 -452
rect -701 -455 -699 -452
rect -692 -455 -690 -452
rect -764 -477 -762 -463
rect -721 -474 -719 -463
rect -764 -484 -762 -481
rect -711 -485 -709 -463
rect -727 -487 -709 -485
rect -764 -507 -762 -504
rect -727 -510 -725 -487
rect -701 -492 -699 -463
rect -711 -494 -699 -492
rect -727 -512 -718 -510
rect -764 -529 -762 -515
rect -720 -529 -718 -512
rect -711 -529 -709 -494
rect -692 -512 -690 -463
rect -702 -514 -690 -512
rect -702 -529 -700 -514
rect -683 -519 -681 -445
rect -58 -455 -56 -452
rect -15 -455 -13 -445
rect -5 -455 -3 -452
rect 5 -455 7 -452
rect 14 -455 16 -452
rect -58 -477 -56 -463
rect -15 -474 -13 -463
rect -58 -484 -56 -481
rect -5 -485 -3 -463
rect -21 -487 -3 -485
rect -58 -507 -56 -504
rect -21 -510 -19 -487
rect 5 -492 7 -463
rect -5 -494 7 -492
rect -21 -512 -12 -510
rect -692 -521 -681 -519
rect -692 -529 -690 -521
rect -58 -529 -56 -515
rect -14 -529 -12 -512
rect -5 -529 -3 -494
rect 14 -512 16 -463
rect 4 -514 16 -512
rect 4 -529 6 -514
rect 23 -519 25 -445
rect 14 -521 25 -519
rect 14 -529 16 -521
rect -764 -536 -762 -533
rect -720 -557 -718 -533
rect -711 -537 -709 -533
rect -702 -568 -700 -533
rect -692 -537 -690 -533
rect -58 -536 -56 -533
rect -14 -557 -12 -533
rect -5 -537 -3 -533
rect 4 -568 6 -533
rect 14 -537 16 -533
rect -714 -693 -712 -690
rect -704 -693 -702 -690
rect -688 -693 -686 -690
rect -536 -693 -534 -690
rect -526 -693 -524 -690
rect -510 -693 -508 -690
rect -356 -693 -354 -690
rect -346 -693 -344 -690
rect -330 -693 -328 -690
rect -145 -693 -143 -690
rect -135 -693 -133 -690
rect -119 -693 -117 -690
rect -714 -725 -712 -701
rect -704 -725 -702 -701
rect -688 -716 -686 -701
rect -714 -732 -712 -729
rect -704 -732 -702 -729
rect -688 -732 -686 -720
rect -536 -725 -534 -701
rect -526 -725 -524 -701
rect -510 -716 -508 -701
rect -536 -732 -534 -729
rect -526 -732 -524 -729
rect -510 -732 -508 -720
rect -356 -725 -354 -701
rect -346 -725 -344 -701
rect -330 -716 -328 -701
rect -356 -732 -354 -729
rect -346 -732 -344 -729
rect -330 -732 -328 -720
rect -145 -725 -143 -701
rect -135 -725 -133 -701
rect -119 -716 -117 -701
rect -145 -732 -143 -729
rect -135 -732 -133 -729
rect -119 -732 -117 -720
rect -785 -838 -783 -828
rect -815 -851 -813 -848
rect -807 -840 -731 -838
rect -807 -851 -805 -840
rect -801 -845 -783 -843
rect -801 -851 -799 -845
rect -793 -851 -791 -848
rect -785 -851 -783 -845
rect -777 -851 -775 -848
rect -771 -851 -769 -840
rect -765 -851 -763 -848
rect -754 -851 -752 -848
rect -741 -851 -739 -848
rect -733 -851 -731 -840
rect -559 -838 -557 -828
rect -725 -851 -723 -848
rect -713 -851 -711 -847
rect -694 -851 -692 -848
rect -589 -851 -587 -848
rect -581 -840 -505 -838
rect -581 -851 -579 -840
rect -575 -845 -557 -843
rect -575 -851 -573 -845
rect -567 -851 -565 -848
rect -559 -851 -557 -845
rect -551 -851 -549 -848
rect -545 -851 -543 -840
rect -539 -851 -537 -848
rect -528 -851 -526 -848
rect -515 -851 -513 -848
rect -507 -851 -505 -840
rect -341 -838 -339 -828
rect -499 -851 -497 -848
rect -487 -851 -485 -847
rect -468 -851 -466 -848
rect -371 -851 -369 -848
rect -363 -840 -287 -838
rect -363 -851 -361 -840
rect -357 -845 -339 -843
rect -357 -851 -355 -845
rect -349 -851 -347 -848
rect -341 -851 -339 -845
rect -333 -851 -331 -848
rect -327 -851 -325 -840
rect -321 -851 -319 -848
rect -310 -851 -308 -848
rect -297 -851 -295 -848
rect -289 -851 -287 -840
rect 18 -845 20 -842
rect 28 -845 30 -842
rect 44 -845 46 -842
rect -281 -851 -279 -848
rect -269 -851 -267 -847
rect -250 -851 -248 -848
rect -815 -861 -813 -859
rect -807 -861 -805 -859
rect -815 -863 -805 -861
rect -815 -902 -813 -863
rect -807 -902 -805 -863
rect -801 -902 -799 -859
rect -793 -902 -791 -859
rect -785 -861 -783 -859
rect -777 -861 -775 -859
rect -785 -863 -775 -861
rect -785 -885 -783 -863
rect -785 -902 -783 -890
rect -777 -902 -775 -863
rect -771 -902 -769 -859
rect -765 -902 -763 -859
rect -754 -894 -752 -859
rect -754 -902 -752 -899
rect -741 -902 -739 -859
rect -733 -902 -731 -859
rect -725 -902 -723 -859
rect -713 -902 -711 -859
rect -694 -902 -692 -859
rect -589 -861 -587 -859
rect -581 -861 -579 -859
rect -589 -863 -579 -861
rect -589 -902 -587 -863
rect -581 -902 -579 -863
rect -575 -902 -573 -859
rect -567 -902 -565 -859
rect -559 -861 -557 -859
rect -551 -861 -549 -859
rect -559 -863 -549 -861
rect -559 -885 -557 -863
rect -559 -902 -557 -890
rect -551 -902 -549 -863
rect -545 -902 -543 -859
rect -539 -902 -537 -859
rect -528 -894 -526 -859
rect -528 -902 -526 -899
rect -515 -902 -513 -859
rect -507 -902 -505 -859
rect -499 -902 -497 -859
rect -487 -902 -485 -859
rect -468 -902 -466 -859
rect -371 -861 -369 -859
rect -363 -861 -361 -859
rect -371 -863 -361 -861
rect -371 -902 -369 -863
rect -363 -902 -361 -863
rect -357 -902 -355 -859
rect -349 -902 -347 -859
rect -341 -861 -339 -859
rect -333 -861 -331 -859
rect -341 -863 -331 -861
rect -341 -885 -339 -863
rect -341 -902 -339 -890
rect -333 -902 -331 -863
rect -327 -902 -325 -859
rect -321 -902 -319 -859
rect -310 -894 -308 -859
rect -310 -902 -308 -899
rect -297 -902 -295 -859
rect -289 -902 -287 -859
rect -281 -902 -279 -859
rect -269 -902 -267 -859
rect -250 -902 -248 -859
rect 18 -877 20 -853
rect 28 -877 30 -853
rect 44 -868 46 -853
rect 18 -884 20 -881
rect 28 -884 30 -881
rect 44 -884 46 -872
rect -825 -911 -822 -907
rect -815 -909 -813 -906
rect -824 -913 -822 -911
rect -807 -909 -805 -906
rect -801 -909 -799 -906
rect -793 -913 -791 -906
rect -785 -909 -783 -906
rect -777 -909 -775 -906
rect -771 -909 -769 -906
rect -765 -913 -763 -906
rect -754 -909 -752 -906
rect -741 -913 -739 -906
rect -733 -909 -731 -906
rect -725 -909 -723 -906
rect -713 -909 -711 -906
rect -694 -909 -692 -906
rect -599 -911 -596 -907
rect -589 -909 -587 -906
rect -824 -915 -812 -913
rect -808 -915 -739 -913
rect -598 -913 -596 -911
rect -581 -909 -579 -906
rect -575 -909 -573 -906
rect -567 -913 -565 -906
rect -559 -909 -557 -906
rect -551 -909 -549 -906
rect -545 -909 -543 -906
rect -539 -913 -537 -906
rect -528 -909 -526 -906
rect -515 -913 -513 -906
rect -507 -909 -505 -906
rect -499 -909 -497 -906
rect -487 -909 -485 -906
rect -468 -909 -466 -906
rect -381 -911 -378 -907
rect -371 -909 -369 -906
rect -598 -915 -586 -913
rect -582 -915 -513 -913
rect -380 -913 -378 -911
rect -363 -909 -361 -906
rect -357 -909 -355 -906
rect -349 -913 -347 -906
rect -341 -909 -339 -906
rect -333 -909 -331 -906
rect -327 -909 -325 -906
rect -321 -913 -319 -906
rect -310 -909 -308 -906
rect -297 -913 -295 -906
rect -289 -909 -287 -906
rect -281 -909 -279 -906
rect -269 -909 -267 -906
rect -250 -909 -248 -906
rect -380 -915 -368 -913
rect -364 -915 -295 -913
rect 4 -915 44 -913
rect -39 -925 -37 -922
rect 4 -925 6 -915
rect 14 -925 16 -922
rect 24 -925 26 -922
rect 33 -925 35 -922
rect -39 -947 -37 -933
rect 4 -944 6 -933
rect -39 -954 -37 -951
rect 14 -955 16 -933
rect -2 -957 16 -955
rect -39 -977 -37 -974
rect -2 -980 0 -957
rect 24 -962 26 -933
rect 14 -964 26 -962
rect -2 -982 7 -980
rect -39 -999 -37 -985
rect 5 -999 7 -982
rect 14 -999 16 -964
rect 33 -982 35 -933
rect 23 -984 35 -982
rect 23 -999 25 -984
rect 42 -989 44 -915
rect 33 -991 44 -989
rect 33 -999 35 -991
rect -39 -1006 -37 -1003
rect 5 -1027 7 -1003
rect 14 -1007 16 -1003
rect 23 -1038 25 -1003
rect 33 -1007 35 -1003
rect -714 -1198 -712 -1195
rect -704 -1198 -702 -1195
rect -688 -1198 -686 -1195
rect -536 -1198 -534 -1195
rect -526 -1198 -524 -1195
rect -510 -1198 -508 -1195
rect -356 -1198 -354 -1195
rect -346 -1198 -344 -1195
rect -330 -1198 -328 -1195
rect -145 -1198 -143 -1195
rect -135 -1198 -133 -1195
rect -119 -1198 -117 -1195
rect -714 -1230 -712 -1206
rect -704 -1230 -702 -1206
rect -688 -1221 -686 -1206
rect -714 -1237 -712 -1234
rect -704 -1237 -702 -1234
rect -688 -1237 -686 -1225
rect -536 -1230 -534 -1206
rect -526 -1230 -524 -1206
rect -510 -1221 -508 -1206
rect -536 -1237 -534 -1234
rect -526 -1237 -524 -1234
rect -510 -1237 -508 -1225
rect -356 -1230 -354 -1206
rect -346 -1230 -344 -1206
rect -330 -1221 -328 -1206
rect -356 -1237 -354 -1234
rect -346 -1237 -344 -1234
rect -330 -1237 -328 -1225
rect -145 -1230 -143 -1206
rect -135 -1230 -133 -1206
rect -119 -1221 -117 -1206
rect -145 -1237 -143 -1234
rect -135 -1237 -133 -1234
rect -119 -1237 -117 -1225
rect -830 -1403 -828 -1393
rect -860 -1416 -858 -1413
rect -852 -1405 -776 -1403
rect -852 -1416 -850 -1405
rect -846 -1410 -828 -1408
rect -846 -1416 -844 -1410
rect -838 -1416 -836 -1413
rect -830 -1416 -828 -1410
rect -822 -1416 -820 -1413
rect -816 -1416 -814 -1405
rect -810 -1416 -808 -1413
rect -799 -1416 -797 -1413
rect -786 -1416 -784 -1413
rect -778 -1416 -776 -1405
rect -604 -1403 -602 -1393
rect -770 -1416 -768 -1413
rect -758 -1416 -756 -1412
rect -739 -1416 -737 -1413
rect -634 -1416 -632 -1413
rect -626 -1405 -550 -1403
rect -626 -1416 -624 -1405
rect -620 -1410 -602 -1408
rect -620 -1416 -618 -1410
rect -612 -1416 -610 -1413
rect -604 -1416 -602 -1410
rect -596 -1416 -594 -1413
rect -590 -1416 -588 -1405
rect -584 -1416 -582 -1413
rect -573 -1416 -571 -1413
rect -560 -1416 -558 -1413
rect -552 -1416 -550 -1405
rect -386 -1403 -384 -1393
rect -544 -1416 -542 -1413
rect -532 -1416 -530 -1412
rect -513 -1416 -511 -1413
rect -416 -1416 -414 -1413
rect -408 -1405 -332 -1403
rect -408 -1416 -406 -1405
rect -402 -1410 -384 -1408
rect -402 -1416 -400 -1410
rect -394 -1416 -392 -1413
rect -386 -1416 -384 -1410
rect -378 -1416 -376 -1413
rect -372 -1416 -370 -1405
rect -366 -1416 -364 -1413
rect -355 -1416 -353 -1413
rect -342 -1416 -340 -1413
rect -334 -1416 -332 -1405
rect 18 -1409 20 -1406
rect 28 -1409 30 -1406
rect 44 -1409 46 -1406
rect -326 -1416 -324 -1413
rect -314 -1416 -312 -1412
rect -295 -1416 -293 -1413
rect -860 -1426 -858 -1424
rect -852 -1426 -850 -1424
rect -860 -1428 -850 -1426
rect -860 -1467 -858 -1428
rect -852 -1467 -850 -1428
rect -846 -1467 -844 -1424
rect -838 -1467 -836 -1424
rect -830 -1426 -828 -1424
rect -822 -1426 -820 -1424
rect -830 -1428 -820 -1426
rect -830 -1450 -828 -1428
rect -830 -1467 -828 -1455
rect -822 -1467 -820 -1428
rect -816 -1467 -814 -1424
rect -810 -1467 -808 -1424
rect -799 -1459 -797 -1424
rect -799 -1467 -797 -1464
rect -786 -1467 -784 -1424
rect -778 -1467 -776 -1424
rect -770 -1467 -768 -1424
rect -758 -1467 -756 -1424
rect -739 -1467 -737 -1424
rect -634 -1426 -632 -1424
rect -626 -1426 -624 -1424
rect -634 -1428 -624 -1426
rect -634 -1467 -632 -1428
rect -626 -1467 -624 -1428
rect -620 -1467 -618 -1424
rect -612 -1467 -610 -1424
rect -604 -1426 -602 -1424
rect -596 -1426 -594 -1424
rect -604 -1428 -594 -1426
rect -604 -1450 -602 -1428
rect -604 -1467 -602 -1455
rect -596 -1467 -594 -1428
rect -590 -1467 -588 -1424
rect -584 -1467 -582 -1424
rect -573 -1459 -571 -1424
rect -573 -1467 -571 -1464
rect -560 -1467 -558 -1424
rect -552 -1467 -550 -1424
rect -544 -1467 -542 -1424
rect -532 -1467 -530 -1424
rect -513 -1467 -511 -1424
rect -416 -1426 -414 -1424
rect -408 -1426 -406 -1424
rect -416 -1428 -406 -1426
rect -416 -1467 -414 -1428
rect -408 -1467 -406 -1428
rect -402 -1467 -400 -1424
rect -394 -1467 -392 -1424
rect -386 -1426 -384 -1424
rect -378 -1426 -376 -1424
rect -386 -1428 -376 -1426
rect -386 -1450 -384 -1428
rect -386 -1467 -384 -1455
rect -378 -1467 -376 -1428
rect -372 -1467 -370 -1424
rect -366 -1467 -364 -1424
rect -355 -1459 -353 -1424
rect -355 -1467 -353 -1464
rect -342 -1467 -340 -1424
rect -334 -1467 -332 -1424
rect -326 -1467 -324 -1424
rect -314 -1467 -312 -1424
rect -295 -1467 -293 -1424
rect 18 -1441 20 -1417
rect 28 -1441 30 -1417
rect 44 -1432 46 -1417
rect 18 -1448 20 -1445
rect 28 -1448 30 -1445
rect 44 -1448 46 -1436
rect -870 -1476 -867 -1472
rect -860 -1474 -858 -1471
rect -869 -1478 -867 -1476
rect -852 -1474 -850 -1471
rect -846 -1474 -844 -1471
rect -838 -1478 -836 -1471
rect -830 -1474 -828 -1471
rect -822 -1474 -820 -1471
rect -816 -1474 -814 -1471
rect -810 -1478 -808 -1471
rect -799 -1474 -797 -1471
rect -786 -1478 -784 -1471
rect -778 -1474 -776 -1471
rect -770 -1474 -768 -1471
rect -758 -1474 -756 -1471
rect -739 -1474 -737 -1471
rect -644 -1476 -641 -1472
rect -634 -1474 -632 -1471
rect -869 -1480 -857 -1478
rect -853 -1480 -784 -1478
rect -643 -1478 -641 -1476
rect -626 -1474 -624 -1471
rect -620 -1474 -618 -1471
rect -612 -1478 -610 -1471
rect -604 -1474 -602 -1471
rect -596 -1474 -594 -1471
rect -590 -1474 -588 -1471
rect -584 -1478 -582 -1471
rect -573 -1474 -571 -1471
rect -560 -1478 -558 -1471
rect -552 -1474 -550 -1471
rect -544 -1474 -542 -1471
rect -532 -1474 -530 -1471
rect -513 -1474 -511 -1471
rect -426 -1476 -423 -1472
rect -416 -1474 -414 -1471
rect -643 -1480 -631 -1478
rect -627 -1480 -558 -1478
rect -425 -1478 -423 -1476
rect -408 -1474 -406 -1471
rect -402 -1474 -400 -1471
rect -394 -1478 -392 -1471
rect -386 -1474 -384 -1471
rect -378 -1474 -376 -1471
rect -372 -1474 -370 -1471
rect -366 -1478 -364 -1471
rect -355 -1474 -353 -1471
rect -342 -1478 -340 -1471
rect -334 -1474 -332 -1471
rect -326 -1474 -324 -1471
rect -314 -1474 -312 -1471
rect -295 -1474 -293 -1471
rect -425 -1480 -413 -1478
rect -409 -1480 -340 -1478
rect 4 -1479 44 -1477
rect -39 -1489 -37 -1486
rect 4 -1489 6 -1479
rect 14 -1489 16 -1486
rect 24 -1489 26 -1486
rect 33 -1489 35 -1486
rect -39 -1511 -37 -1497
rect 4 -1508 6 -1497
rect -39 -1518 -37 -1515
rect 14 -1519 16 -1497
rect -2 -1521 16 -1519
rect -39 -1541 -37 -1538
rect -2 -1544 0 -1521
rect 24 -1526 26 -1497
rect 14 -1528 26 -1526
rect -2 -1546 7 -1544
rect -39 -1563 -37 -1549
rect 5 -1563 7 -1546
rect 14 -1563 16 -1528
rect 33 -1546 35 -1497
rect 23 -1548 35 -1546
rect 23 -1563 25 -1548
rect 42 -1553 44 -1479
rect 33 -1555 44 -1553
rect 33 -1563 35 -1555
rect -39 -1570 -37 -1567
rect 5 -1591 7 -1567
rect 14 -1571 16 -1567
rect 23 -1602 25 -1567
rect 33 -1571 35 -1567
<< polycontact >>
rect -333 -9 -329 -5
rect -323 -17 -319 -13
rect -307 -9 -303 -5
rect -212 -9 -208 -5
rect -202 -17 -198 -13
rect -186 -9 -182 -5
rect -98 -9 -94 -5
rect -88 -17 -84 -13
rect -72 -9 -68 -5
rect 2 -9 6 -5
rect 12 -17 16 -13
rect 28 -9 32 -5
rect -433 -227 -429 -223
rect -423 -235 -419 -231
rect -407 -227 -403 -223
rect -275 -227 -271 -223
rect -265 -235 -261 -231
rect -249 -227 -245 -223
rect -136 -227 -132 -223
rect -126 -235 -122 -231
rect -110 -227 -106 -223
rect -18 -227 -14 -223
rect -8 -235 -4 -231
rect 8 -227 12 -223
rect -564 -358 -560 -354
rect -312 -358 -308 -354
rect -711 -395 -707 -391
rect -701 -403 -697 -399
rect -685 -395 -681 -391
rect -495 -409 -491 -405
rect -243 -409 -239 -405
rect -5 -395 -1 -391
rect 5 -403 9 -399
rect 21 -395 25 -391
rect -606 -441 -602 -437
rect -354 -442 -350 -438
rect -768 -474 -764 -470
rect -725 -474 -721 -470
rect -715 -497 -711 -493
rect -768 -526 -764 -522
rect -62 -474 -58 -470
rect -19 -474 -15 -470
rect -9 -497 -5 -493
rect -62 -526 -58 -522
rect -724 -557 -720 -553
rect -706 -568 -702 -564
rect -18 -557 -14 -553
rect 0 -568 4 -564
rect -718 -713 -714 -709
rect -708 -721 -704 -717
rect -692 -713 -688 -709
rect -540 -713 -536 -709
rect -530 -721 -526 -717
rect -514 -713 -510 -709
rect -360 -713 -356 -709
rect -350 -721 -346 -717
rect -334 -713 -330 -709
rect -149 -713 -145 -709
rect -139 -721 -135 -717
rect -123 -713 -119 -709
rect -786 -828 -782 -824
rect -560 -828 -556 -824
rect -342 -828 -338 -824
rect -717 -879 -713 -875
rect -491 -879 -487 -875
rect -273 -879 -269 -875
rect 14 -865 18 -861
rect 24 -873 28 -869
rect 40 -865 44 -861
rect -829 -911 -825 -907
rect -603 -911 -599 -907
rect -385 -911 -381 -907
rect -43 -944 -39 -940
rect 0 -944 4 -940
rect 10 -967 14 -963
rect -43 -996 -39 -992
rect 1 -1027 5 -1023
rect 19 -1038 23 -1034
rect -718 -1218 -714 -1214
rect -708 -1226 -704 -1222
rect -692 -1218 -688 -1214
rect -540 -1218 -536 -1214
rect -530 -1226 -526 -1222
rect -514 -1218 -510 -1214
rect -360 -1218 -356 -1214
rect -350 -1226 -346 -1222
rect -334 -1218 -330 -1214
rect -149 -1218 -145 -1214
rect -139 -1226 -135 -1222
rect -123 -1218 -119 -1214
rect -831 -1393 -827 -1389
rect -605 -1393 -601 -1389
rect -387 -1393 -383 -1389
rect -762 -1444 -758 -1440
rect -536 -1444 -532 -1440
rect -318 -1444 -314 -1440
rect 14 -1429 18 -1425
rect 24 -1437 28 -1433
rect 40 -1429 44 -1425
rect -874 -1476 -870 -1472
rect -648 -1476 -644 -1472
rect -430 -1476 -426 -1472
rect -43 -1508 -39 -1504
rect 0 -1508 4 -1504
rect 10 -1531 14 -1527
rect -43 -1560 -39 -1556
rect 1 -1591 5 -1587
rect 19 -1602 23 -1598
<< metal1 >>
rect -345 101 273 106
rect -223 79 217 84
rect -109 58 159 63
rect -9 36 118 42
rect -951 17 45 21
rect -995 -247 -991 -33
rect -951 -197 -947 17
rect -334 11 -330 17
rect -316 11 -312 17
rect -308 11 -304 17
rect -213 11 -209 17
rect -195 11 -191 17
rect -187 11 -183 17
rect -99 11 -95 17
rect -81 11 -77 17
rect -73 11 -69 17
rect 1 11 5 17
rect 19 11 23 17
rect 27 11 31 17
rect -324 0 -320 3
rect -324 -3 -312 0
rect -316 -5 -312 -3
rect -300 -5 -296 3
rect -203 0 -199 3
rect -203 -3 -191 0
rect -345 -9 -333 -5
rect -316 -9 -307 -5
rect -300 -9 -283 -5
rect -195 -5 -191 -3
rect -179 -5 -175 3
rect -89 0 -85 3
rect -89 -3 -77 0
rect -223 -9 -212 -5
rect -195 -9 -186 -5
rect -179 -9 -159 -5
rect -81 -5 -77 -3
rect -65 -5 -61 3
rect 11 0 15 3
rect 11 -3 23 0
rect -109 -9 -98 -5
rect -81 -9 -72 -5
rect -65 -9 -49 -5
rect 19 -5 23 -3
rect 35 -5 39 3
rect -9 -9 2 -5
rect 19 -9 28 -5
rect 35 -9 64 -5
rect -359 -17 -323 -13
rect -316 -21 -312 -9
rect -300 -12 -296 -9
rect -334 -29 -330 -25
rect -308 -29 -304 -16
rect -237 -17 -202 -13
rect -195 -21 -191 -9
rect -179 -12 -175 -9
rect -213 -29 -209 -25
rect -187 -29 -183 -16
rect -123 -17 -88 -13
rect -81 -21 -77 -9
rect -65 -12 -61 -9
rect -99 -29 -95 -25
rect -73 -29 -69 -16
rect -23 -17 12 -13
rect 19 -21 23 -9
rect 35 -12 39 -9
rect 1 -29 5 -25
rect 27 -29 31 -16
rect -919 -33 45 -29
rect -332 -46 -159 -42
rect -74 -46 -49 -42
rect -332 -87 -328 -46
rect -74 -91 -70 -46
rect -444 -118 63 -113
rect -286 -139 65 -134
rect -147 -158 58 -153
rect 63 -158 64 -153
rect 95 -176 101 36
rect 100 -181 101 -176
rect -951 -201 25 -197
rect -995 -251 -965 -247
rect -995 -543 -991 -251
rect -951 -367 -947 -201
rect -434 -207 -430 -201
rect -416 -207 -412 -201
rect -408 -207 -404 -201
rect -276 -207 -272 -201
rect -258 -207 -254 -201
rect -250 -207 -246 -201
rect -137 -207 -133 -201
rect -119 -207 -115 -201
rect -111 -207 -107 -201
rect -19 -207 -15 -201
rect -1 -207 3 -201
rect 7 -207 11 -201
rect -424 -218 -420 -215
rect -424 -221 -412 -218
rect -416 -223 -412 -221
rect -400 -223 -396 -215
rect -266 -218 -262 -215
rect -266 -221 -254 -218
rect -444 -227 -433 -223
rect -416 -227 -407 -223
rect -400 -227 -379 -223
rect -258 -223 -254 -221
rect -242 -223 -238 -215
rect -127 -218 -123 -215
rect -127 -221 -115 -218
rect -286 -227 -275 -223
rect -258 -227 -249 -223
rect -242 -227 -232 -223
rect -119 -223 -115 -221
rect -103 -223 -99 -215
rect -9 -218 -5 -215
rect -9 -221 3 -218
rect -147 -227 -136 -223
rect -119 -227 -110 -223
rect -103 -227 -92 -223
rect -1 -223 3 -221
rect 15 -223 19 -215
rect -29 -227 -18 -223
rect -1 -227 8 -223
rect 15 -227 56 -223
rect -458 -235 -423 -231
rect -416 -239 -412 -227
rect -400 -230 -396 -227
rect -434 -247 -430 -243
rect -408 -247 -404 -234
rect -300 -235 -265 -231
rect -258 -239 -254 -227
rect -242 -230 -238 -227
rect -276 -247 -272 -243
rect -250 -247 -246 -234
rect -161 -235 -126 -231
rect -119 -239 -115 -227
rect -103 -230 -99 -227
rect -137 -247 -133 -243
rect -111 -247 -107 -234
rect -43 -235 -8 -231
rect -1 -239 3 -227
rect 15 -230 19 -227
rect -19 -247 -15 -243
rect 7 -247 11 -234
rect -926 -251 25 -247
rect -571 -275 -538 -271
rect -861 -336 -646 -332
rect -564 -354 -560 -307
rect -332 -354 -328 -288
rect -332 -358 -312 -354
rect -811 -367 -590 -366
rect -951 -369 -590 -367
rect -951 -371 -807 -369
rect -995 -547 -977 -543
rect -995 -733 -991 -547
rect -951 -683 -947 -371
rect -811 -445 -807 -371
rect -712 -375 -708 -369
rect -694 -375 -690 -369
rect -686 -375 -682 -369
rect -604 -370 -590 -369
rect -586 -370 -338 -366
rect -334 -369 38 -366
rect -334 -370 -101 -369
rect -702 -386 -698 -383
rect -702 -389 -690 -386
rect -694 -391 -690 -389
rect -678 -391 -674 -383
rect -598 -377 -564 -373
rect -598 -381 -594 -377
rect -568 -381 -564 -377
rect -560 -381 -556 -370
rect -516 -381 -512 -370
rect -498 -381 -494 -370
rect -477 -381 -473 -370
rect -346 -377 -312 -373
rect -346 -381 -342 -377
rect -316 -381 -312 -377
rect -799 -395 -711 -391
rect -694 -395 -685 -391
rect -678 -395 -646 -391
rect -790 -403 -701 -399
rect -694 -407 -690 -395
rect -678 -398 -674 -395
rect -712 -415 -708 -411
rect -686 -415 -682 -402
rect -718 -419 -672 -415
rect -576 -424 -572 -389
rect -540 -405 -536 -389
rect -308 -381 -304 -370
rect -264 -381 -260 -370
rect -246 -381 -242 -370
rect -225 -381 -221 -370
rect -526 -392 -522 -389
rect -508 -392 -504 -389
rect -526 -396 -504 -392
rect -486 -401 -482 -389
rect -540 -409 -495 -405
rect -540 -416 -536 -409
rect -522 -420 -504 -416
rect -576 -428 -532 -424
rect -576 -432 -572 -428
rect -508 -432 -504 -420
rect -486 -432 -482 -406
rect -469 -413 -465 -389
rect -456 -405 -411 -401
rect -469 -417 -446 -413
rect -469 -432 -465 -417
rect -324 -424 -320 -389
rect -288 -405 -284 -389
rect -274 -392 -270 -389
rect -256 -392 -252 -389
rect -274 -396 -252 -392
rect -234 -401 -230 -389
rect -288 -409 -243 -405
rect -288 -416 -284 -409
rect -270 -420 -252 -416
rect -324 -428 -280 -424
rect -324 -432 -320 -428
rect -256 -432 -252 -420
rect -234 -432 -230 -406
rect -217 -413 -213 -389
rect -204 -405 -190 -401
rect -217 -417 -204 -413
rect -217 -432 -213 -417
rect -618 -441 -606 -437
rect -598 -441 -594 -436
rect -568 -441 -564 -436
rect -598 -445 -564 -441
rect -811 -449 -675 -445
rect -560 -449 -556 -436
rect -516 -449 -512 -436
rect -498 -449 -494 -436
rect -477 -449 -473 -436
rect -362 -442 -354 -438
rect -346 -441 -342 -436
rect -316 -441 -312 -436
rect -346 -445 -312 -441
rect -308 -449 -304 -436
rect -264 -449 -260 -436
rect -246 -449 -242 -436
rect -225 -449 -221 -436
rect -105 -445 -101 -370
rect -6 -375 -2 -369
rect 12 -375 16 -369
rect 20 -375 24 -369
rect 4 -386 8 -383
rect 4 -389 16 -386
rect 12 -391 16 -389
rect 28 -391 32 -383
rect -93 -395 -5 -391
rect 12 -395 21 -391
rect 28 -395 62 -391
rect -84 -403 5 -399
rect 12 -407 16 -395
rect 28 -398 32 -395
rect -6 -415 -2 -411
rect 20 -415 24 -402
rect -12 -419 34 -415
rect -105 -449 33 -445
rect -841 -489 -796 -485
rect -784 -497 -780 -449
rect -769 -455 -765 -449
rect -727 -455 -723 -449
rect -689 -455 -685 -449
rect -645 -453 -590 -449
rect -586 -453 -338 -449
rect -334 -453 -155 -449
rect -761 -470 -757 -463
rect -772 -474 -768 -470
rect -761 -474 -725 -470
rect -761 -477 -757 -474
rect -769 -487 -765 -481
rect -772 -491 -744 -487
rect -784 -501 -751 -497
rect -769 -507 -765 -501
rect -748 -510 -744 -491
rect -735 -497 -715 -493
rect -707 -501 -703 -463
rect -707 -505 -663 -501
rect -748 -514 -734 -510
rect -838 -526 -812 -522
rect -761 -522 -757 -515
rect -806 -526 -797 -522
rect -893 -547 -851 -543
rect -838 -573 -834 -526
rect -792 -526 -768 -522
rect -761 -526 -754 -522
rect -761 -529 -757 -526
rect -769 -543 -765 -533
rect -738 -543 -734 -514
rect -707 -529 -703 -505
rect -727 -543 -723 -533
rect -689 -543 -685 -533
rect -805 -547 -672 -543
rect -689 -552 -685 -547
rect -645 -552 -641 -453
rect -790 -557 -724 -553
rect -689 -556 -641 -552
rect -747 -568 -706 -564
rect -446 -573 -442 -464
rect -838 -577 -442 -573
rect -639 -609 -635 -591
rect -411 -610 -407 -461
rect -362 -474 -176 -470
rect -190 -606 -186 -575
rect -180 -585 -176 -474
rect -159 -543 -155 -453
rect -122 -474 -91 -470
rect -78 -497 -74 -449
rect -63 -455 -59 -449
rect -21 -455 -17 -449
rect 17 -455 21 -449
rect -55 -470 -51 -463
rect -66 -474 -62 -470
rect -55 -474 -19 -470
rect -55 -477 -51 -474
rect -63 -487 -59 -481
rect -66 -491 -38 -487
rect -78 -501 -45 -497
rect -63 -507 -59 -501
rect -42 -510 -38 -491
rect -29 -497 -9 -493
rect -1 -501 3 -463
rect -1 -505 45 -501
rect -42 -514 -28 -510
rect -138 -526 -106 -522
rect -55 -522 -51 -515
rect -100 -526 -91 -522
rect -86 -526 -62 -522
rect -55 -526 -48 -522
rect -55 -529 -51 -526
rect -63 -543 -59 -533
rect -32 -543 -28 -514
rect -1 -529 3 -505
rect -21 -543 -17 -533
rect 17 -543 21 -533
rect -159 -547 34 -543
rect -84 -557 -18 -553
rect -41 -568 0 -564
rect 58 -585 62 -395
rect -180 -589 62 -585
rect -729 -624 42 -619
rect -551 -639 40 -634
rect 45 -639 47 -634
rect -372 -659 -7 -654
rect 95 -670 101 -181
rect -160 -675 94 -670
rect -951 -687 -91 -683
rect -997 -737 -970 -733
rect -995 -919 -991 -737
rect -951 -836 -947 -687
rect -719 -693 -715 -687
rect -701 -693 -697 -687
rect -693 -693 -689 -687
rect -541 -693 -537 -687
rect -523 -693 -519 -687
rect -515 -693 -511 -687
rect -361 -693 -357 -687
rect -343 -693 -339 -687
rect -335 -693 -331 -687
rect -150 -693 -146 -687
rect -132 -693 -128 -687
rect -124 -693 -120 -687
rect -709 -704 -705 -701
rect -709 -707 -697 -704
rect -701 -709 -697 -707
rect -685 -709 -681 -701
rect -531 -704 -527 -701
rect -531 -707 -519 -704
rect -729 -713 -718 -709
rect -701 -713 -692 -709
rect -685 -713 -675 -709
rect -523 -709 -519 -707
rect -507 -709 -503 -701
rect -351 -704 -347 -701
rect -351 -707 -339 -704
rect -551 -713 -540 -709
rect -523 -713 -514 -709
rect -507 -713 -497 -709
rect -343 -709 -339 -707
rect -327 -709 -323 -701
rect -140 -704 -136 -701
rect -140 -707 -128 -704
rect -371 -713 -360 -709
rect -343 -713 -334 -709
rect -327 -713 -317 -709
rect -132 -709 -128 -707
rect -116 -709 -112 -701
rect -160 -713 -149 -709
rect -132 -713 -123 -709
rect -116 -713 -106 -709
rect -743 -721 -708 -717
rect -701 -725 -697 -713
rect -685 -716 -681 -713
rect -719 -733 -715 -729
rect -693 -733 -689 -720
rect -565 -721 -530 -717
rect -523 -725 -519 -713
rect -507 -716 -503 -713
rect -541 -733 -537 -729
rect -515 -733 -511 -720
rect -385 -721 -350 -717
rect -343 -725 -339 -713
rect -327 -716 -323 -713
rect -361 -733 -357 -729
rect -335 -733 -331 -720
rect -174 -721 -139 -717
rect -132 -725 -128 -713
rect -116 -716 -112 -713
rect -150 -733 -146 -729
rect -124 -733 -120 -720
rect -904 -737 -91 -733
rect -861 -791 -782 -787
rect -786 -824 -782 -791
rect -406 -800 -338 -796
rect -561 -823 -557 -807
rect -560 -824 -556 -823
rect -342 -824 -338 -800
rect -951 -840 -812 -836
rect -808 -840 -586 -836
rect -582 -840 -368 -836
rect -364 -839 57 -836
rect -364 -840 -82 -839
rect -996 -923 -974 -919
rect -995 -1238 -991 -923
rect -951 -1188 -947 -840
rect -820 -847 -786 -843
rect -820 -851 -816 -847
rect -790 -851 -786 -847
rect -782 -851 -778 -840
rect -738 -851 -734 -840
rect -720 -851 -716 -840
rect -699 -851 -695 -840
rect -594 -847 -560 -843
rect -594 -851 -590 -847
rect -564 -851 -560 -847
rect -798 -894 -794 -859
rect -762 -875 -758 -859
rect -556 -851 -552 -840
rect -512 -851 -508 -840
rect -494 -851 -490 -840
rect -473 -851 -469 -840
rect -376 -847 -342 -843
rect -376 -851 -372 -847
rect -346 -851 -342 -847
rect -748 -862 -744 -859
rect -730 -862 -726 -859
rect -748 -866 -726 -862
rect -708 -871 -704 -859
rect -762 -879 -717 -875
rect -762 -886 -758 -879
rect -744 -890 -726 -886
rect -798 -898 -754 -894
rect -798 -902 -794 -898
rect -730 -902 -726 -890
rect -708 -902 -704 -876
rect -691 -883 -687 -859
rect -678 -875 -661 -871
rect -691 -887 -678 -883
rect -691 -902 -687 -887
rect -572 -894 -568 -859
rect -536 -875 -532 -859
rect -338 -851 -334 -840
rect -294 -851 -290 -840
rect -276 -851 -272 -840
rect -255 -851 -251 -840
rect -522 -862 -518 -859
rect -504 -862 -500 -859
rect -522 -866 -500 -862
rect -482 -871 -478 -859
rect -536 -879 -491 -875
rect -536 -886 -532 -879
rect -518 -890 -500 -886
rect -572 -898 -528 -894
rect -572 -902 -568 -898
rect -504 -902 -500 -890
rect -482 -902 -478 -876
rect -465 -883 -461 -859
rect -452 -875 -422 -871
rect -465 -887 -447 -883
rect -465 -902 -461 -887
rect -354 -894 -350 -859
rect -318 -875 -314 -859
rect -304 -862 -300 -859
rect -286 -862 -282 -859
rect -304 -866 -282 -862
rect -264 -871 -260 -859
rect -318 -879 -273 -875
rect -318 -886 -314 -879
rect -300 -890 -282 -886
rect -354 -898 -310 -894
rect -354 -902 -350 -898
rect -286 -902 -282 -890
rect -264 -902 -260 -876
rect -247 -883 -243 -859
rect -234 -875 -203 -871
rect -247 -887 -221 -883
rect -247 -902 -243 -887
rect -844 -911 -829 -907
rect -820 -911 -816 -906
rect -790 -911 -786 -906
rect -844 -946 -840 -911
rect -820 -915 -786 -911
rect -782 -919 -778 -906
rect -738 -919 -734 -906
rect -720 -919 -716 -906
rect -699 -919 -695 -906
rect -614 -911 -603 -907
rect -594 -911 -590 -906
rect -564 -911 -560 -906
rect -594 -915 -560 -911
rect -556 -919 -552 -906
rect -512 -919 -508 -906
rect -494 -919 -490 -906
rect -473 -919 -469 -906
rect -396 -911 -385 -907
rect -376 -911 -372 -906
rect -346 -911 -342 -906
rect -376 -915 -342 -911
rect -338 -919 -334 -906
rect -294 -919 -290 -906
rect -276 -919 -272 -906
rect -255 -919 -251 -906
rect -826 -923 -812 -919
rect -808 -923 -586 -919
rect -582 -923 -368 -919
rect -364 -923 -235 -919
rect -844 -950 -447 -946
rect -660 -1109 -656 -1081
rect -422 -1109 -418 -944
rect -396 -947 -252 -943
rect -256 -1049 -252 -947
rect -239 -1013 -235 -923
rect -225 -973 -221 -887
rect -207 -991 -203 -875
rect -86 -915 -82 -840
rect 13 -845 17 -839
rect 31 -845 35 -839
rect 39 -845 43 -839
rect 23 -856 27 -853
rect 23 -859 35 -856
rect 31 -861 35 -859
rect 47 -861 51 -853
rect -74 -865 14 -861
rect 31 -865 40 -861
rect 47 -865 77 -861
rect -65 -873 24 -869
rect 31 -877 35 -865
rect 47 -868 51 -865
rect 13 -885 17 -881
rect 39 -885 43 -872
rect 7 -889 53 -885
rect -86 -919 50 -915
rect -101 -944 -72 -940
rect -59 -967 -55 -919
rect -44 -925 -40 -919
rect -2 -925 2 -919
rect 36 -925 40 -919
rect -36 -940 -32 -933
rect -47 -944 -43 -940
rect -36 -944 0 -940
rect -36 -947 -32 -944
rect -44 -957 -40 -951
rect -47 -961 -19 -957
rect -59 -971 -26 -967
rect -44 -977 -40 -971
rect -23 -980 -19 -961
rect -10 -967 10 -963
rect 18 -971 22 -933
rect 18 -975 62 -971
rect -23 -984 -9 -980
rect -185 -996 -87 -992
rect -36 -992 -32 -985
rect -81 -996 -72 -992
rect -67 -996 -43 -992
rect -36 -996 -29 -992
rect -36 -999 -32 -996
rect -44 -1013 -40 -1003
rect -13 -1013 -9 -984
rect 18 -999 22 -975
rect -2 -1013 2 -1003
rect 36 -1013 40 -1003
rect -239 -1017 53 -1013
rect -65 -1027 1 -1023
rect -22 -1038 19 -1034
rect 73 -1049 77 -865
rect -256 -1053 77 -1049
rect -207 -1110 -203 -1070
rect -729 -1129 42 -1124
rect -551 -1144 40 -1139
rect 45 -1144 47 -1139
rect -372 -1164 -7 -1159
rect 84 -1166 88 -1089
rect 95 -1175 101 -675
rect 141 -153 146 58
rect 141 -654 146 -158
rect 141 -1159 146 -659
rect 187 -134 192 79
rect 187 -634 192 -139
rect 187 -1139 192 -639
rect 247 -113 252 101
rect 308 -80 371 -76
rect 247 -619 252 -118
rect 247 -624 248 -619
rect 247 -1124 252 -624
rect 285 -676 289 -505
rect 331 -634 335 -568
rect 264 -1105 299 -1101
rect 331 -1119 335 -1068
rect 247 -1129 248 -1124
rect -160 -1180 94 -1175
rect -951 -1192 -91 -1188
rect -996 -1242 -974 -1238
rect -995 -1484 -991 -1242
rect -951 -1401 -947 -1192
rect -719 -1198 -715 -1192
rect -701 -1198 -697 -1192
rect -693 -1198 -689 -1192
rect -541 -1198 -537 -1192
rect -523 -1198 -519 -1192
rect -515 -1198 -511 -1192
rect -361 -1198 -357 -1192
rect -343 -1198 -339 -1192
rect -335 -1198 -331 -1192
rect -150 -1198 -146 -1192
rect -132 -1198 -128 -1192
rect -124 -1198 -120 -1192
rect -709 -1209 -705 -1206
rect -709 -1212 -697 -1209
rect -701 -1214 -697 -1212
rect -685 -1214 -681 -1206
rect -531 -1209 -527 -1206
rect -531 -1212 -519 -1209
rect -729 -1218 -718 -1214
rect -701 -1218 -692 -1214
rect -685 -1218 -675 -1214
rect -523 -1214 -519 -1212
rect -507 -1214 -503 -1206
rect -351 -1209 -347 -1206
rect -351 -1212 -339 -1209
rect -551 -1218 -540 -1214
rect -523 -1218 -514 -1214
rect -507 -1218 -497 -1214
rect -343 -1214 -339 -1212
rect -327 -1214 -323 -1206
rect -140 -1209 -136 -1206
rect -140 -1212 -128 -1209
rect -371 -1218 -360 -1214
rect -343 -1218 -334 -1214
rect -327 -1218 -317 -1214
rect -132 -1214 -128 -1212
rect -116 -1214 -112 -1206
rect -160 -1218 -149 -1214
rect -132 -1218 -123 -1214
rect -116 -1218 -106 -1214
rect -743 -1226 -708 -1222
rect -701 -1230 -697 -1218
rect -685 -1221 -681 -1218
rect -719 -1238 -715 -1234
rect -693 -1238 -689 -1225
rect -565 -1226 -530 -1222
rect -523 -1230 -519 -1218
rect -507 -1221 -503 -1218
rect -541 -1238 -537 -1234
rect -515 -1238 -511 -1225
rect -385 -1226 -350 -1222
rect -343 -1230 -339 -1218
rect -327 -1221 -323 -1218
rect -361 -1238 -357 -1234
rect -335 -1238 -331 -1225
rect -174 -1226 -139 -1222
rect -132 -1230 -128 -1218
rect -116 -1221 -112 -1218
rect -150 -1238 -146 -1234
rect -124 -1238 -120 -1225
rect -915 -1242 -91 -1238
rect -656 -1318 -601 -1314
rect -831 -1389 -827 -1350
rect -605 -1389 -601 -1318
rect -418 -1337 -383 -1333
rect -387 -1389 -383 -1337
rect -257 -1401 57 -1400
rect -952 -1405 -857 -1401
rect -853 -1405 -631 -1401
rect -627 -1405 -413 -1401
rect -409 -1403 57 -1401
rect -409 -1404 -82 -1403
rect -409 -1405 -251 -1404
rect -865 -1412 -831 -1408
rect -865 -1416 -861 -1412
rect -835 -1416 -831 -1412
rect -827 -1416 -823 -1405
rect -783 -1416 -779 -1405
rect -765 -1416 -761 -1405
rect -744 -1416 -740 -1405
rect -639 -1412 -605 -1408
rect -639 -1416 -635 -1412
rect -609 -1416 -605 -1412
rect -843 -1459 -839 -1424
rect -807 -1440 -803 -1424
rect -601 -1416 -597 -1405
rect -557 -1416 -553 -1405
rect -539 -1416 -535 -1405
rect -518 -1416 -514 -1405
rect -421 -1412 -387 -1408
rect -421 -1416 -417 -1412
rect -391 -1416 -387 -1412
rect -793 -1427 -789 -1424
rect -775 -1427 -771 -1424
rect -793 -1431 -771 -1427
rect -753 -1436 -749 -1424
rect -807 -1444 -762 -1440
rect -807 -1451 -803 -1444
rect -789 -1455 -771 -1451
rect -843 -1463 -799 -1459
rect -843 -1467 -839 -1463
rect -775 -1467 -771 -1455
rect -753 -1467 -749 -1441
rect -736 -1448 -732 -1424
rect -723 -1440 -693 -1436
rect -736 -1452 -724 -1448
rect -736 -1467 -732 -1452
rect -617 -1459 -613 -1424
rect -581 -1440 -577 -1424
rect -383 -1416 -379 -1405
rect -339 -1416 -335 -1405
rect -321 -1416 -317 -1405
rect -300 -1416 -296 -1405
rect -567 -1427 -563 -1424
rect -549 -1427 -545 -1424
rect -567 -1431 -545 -1427
rect -527 -1436 -523 -1424
rect -581 -1444 -536 -1440
rect -581 -1451 -577 -1444
rect -563 -1455 -545 -1451
rect -617 -1463 -573 -1459
rect -617 -1467 -613 -1463
rect -549 -1467 -545 -1455
rect -527 -1467 -523 -1441
rect -510 -1448 -506 -1424
rect -497 -1440 -469 -1436
rect -510 -1452 -492 -1448
rect -510 -1467 -506 -1452
rect -399 -1459 -395 -1424
rect -363 -1440 -359 -1424
rect -349 -1427 -345 -1424
rect -331 -1427 -327 -1424
rect -349 -1431 -327 -1427
rect -309 -1436 -305 -1424
rect -363 -1444 -318 -1440
rect -363 -1451 -359 -1444
rect -345 -1455 -327 -1451
rect -399 -1463 -355 -1459
rect -399 -1467 -395 -1463
rect -331 -1467 -327 -1455
rect -309 -1467 -305 -1441
rect -292 -1448 -288 -1424
rect -279 -1440 -242 -1436
rect -292 -1452 -266 -1448
rect -292 -1467 -288 -1452
rect -888 -1476 -874 -1472
rect -865 -1476 -861 -1471
rect -835 -1476 -831 -1471
rect -865 -1480 -831 -1476
rect -827 -1484 -823 -1471
rect -783 -1484 -779 -1471
rect -765 -1484 -761 -1471
rect -744 -1484 -740 -1471
rect -659 -1476 -648 -1472
rect -639 -1476 -635 -1471
rect -609 -1476 -605 -1471
rect -639 -1480 -605 -1476
rect -601 -1484 -597 -1471
rect -557 -1484 -553 -1471
rect -539 -1484 -535 -1471
rect -518 -1484 -514 -1471
rect -441 -1476 -430 -1472
rect -421 -1476 -417 -1471
rect -391 -1476 -387 -1471
rect -421 -1480 -387 -1476
rect -383 -1484 -379 -1471
rect -339 -1484 -335 -1471
rect -321 -1484 -317 -1471
rect -300 -1484 -296 -1471
rect -996 -1488 -857 -1484
rect -853 -1488 -631 -1484
rect -627 -1488 -413 -1484
rect -409 -1488 -280 -1484
rect -724 -1699 -720 -1513
rect -640 -1510 -423 -1506
rect -693 -1699 -689 -1513
rect -284 -1577 -280 -1488
rect -270 -1505 -266 -1452
rect -86 -1479 -82 -1404
rect 13 -1409 17 -1403
rect 31 -1409 35 -1403
rect 39 -1409 43 -1403
rect 23 -1420 27 -1417
rect 23 -1423 35 -1420
rect 31 -1425 35 -1423
rect 47 -1425 51 -1417
rect -74 -1429 14 -1425
rect 31 -1429 40 -1425
rect 47 -1429 77 -1425
rect -65 -1437 24 -1433
rect 31 -1441 35 -1429
rect 47 -1432 51 -1429
rect 13 -1449 17 -1445
rect 39 -1449 43 -1436
rect 7 -1453 53 -1449
rect -86 -1483 50 -1479
rect -101 -1508 -72 -1504
rect -59 -1531 -55 -1483
rect -44 -1489 -40 -1483
rect -2 -1489 2 -1483
rect 36 -1489 40 -1483
rect -36 -1504 -32 -1497
rect -47 -1508 -43 -1504
rect -36 -1508 0 -1504
rect -36 -1511 -32 -1508
rect -44 -1521 -40 -1515
rect -47 -1525 -19 -1521
rect -59 -1535 -26 -1531
rect -44 -1541 -40 -1535
rect -23 -1544 -19 -1525
rect -10 -1531 10 -1527
rect 18 -1535 22 -1497
rect 18 -1539 62 -1535
rect -23 -1548 -9 -1544
rect -202 -1560 -87 -1556
rect -36 -1556 -32 -1549
rect -81 -1560 -72 -1556
rect -67 -1560 -43 -1556
rect -36 -1560 -29 -1556
rect -36 -1563 -32 -1560
rect -44 -1577 -40 -1567
rect -13 -1577 -9 -1548
rect 18 -1563 22 -1539
rect -2 -1577 2 -1567
rect 36 -1577 40 -1567
rect -284 -1581 53 -1577
rect -65 -1591 1 -1587
rect -22 -1602 19 -1598
rect 73 -1613 77 -1429
rect -442 -1617 77 -1613
<< m2contact >>
rect -350 101 -345 106
rect -228 79 -223 84
rect -114 58 -109 63
rect -15 36 -9 42
rect -995 -33 -990 -28
rect -350 -9 -345 -4
rect -283 -9 -278 -4
rect -228 -9 -223 -4
rect -159 -9 -154 -4
rect -114 -9 -109 -4
rect -49 -9 -44 -4
rect -14 -9 -9 -4
rect 64 -9 69 -4
rect -364 -17 -359 -12
rect -242 -17 -237 -12
rect -128 -17 -123 -12
rect -28 -17 -23 -12
rect -923 -33 -919 -29
rect -159 -46 -154 -41
rect -49 -46 -44 -41
rect -332 -92 -327 -87
rect -74 -95 -70 -91
rect -449 -118 -444 -113
rect 63 -118 68 -113
rect -291 -139 -286 -134
rect 65 -139 70 -134
rect -152 -158 -147 -153
rect 58 -158 63 -153
rect 95 -181 100 -176
rect -965 -251 -960 -246
rect -449 -227 -444 -222
rect -379 -227 -374 -222
rect -291 -227 -286 -222
rect -232 -227 -227 -222
rect -152 -227 -147 -222
rect -92 -227 -88 -223
rect -34 -227 -29 -222
rect 56 -227 61 -222
rect -463 -235 -458 -230
rect -931 -251 -926 -246
rect -305 -235 -300 -230
rect -166 -235 -161 -230
rect -48 -235 -43 -230
rect -576 -275 -571 -270
rect -538 -275 -533 -270
rect -332 -288 -327 -283
rect -564 -307 -559 -302
rect -866 -336 -861 -331
rect -646 -336 -641 -331
rect -977 -547 -972 -542
rect -804 -396 -799 -391
rect -646 -395 -641 -390
rect -795 -404 -790 -399
rect -672 -419 -667 -414
rect -486 -406 -481 -401
rect -461 -406 -456 -401
rect -411 -405 -406 -400
rect -446 -417 -441 -412
rect -234 -406 -229 -401
rect -209 -406 -204 -401
rect -190 -405 -185 -400
rect -204 -417 -199 -412
rect -624 -441 -618 -435
rect -367 -442 -362 -437
rect -98 -396 -93 -391
rect -89 -404 -84 -399
rect 34 -419 39 -414
rect -846 -490 -841 -485
rect -796 -489 -791 -484
rect -777 -475 -772 -470
rect -740 -498 -735 -493
rect -663 -505 -658 -500
rect -812 -526 -806 -520
rect -898 -547 -893 -542
rect -851 -547 -846 -542
rect -797 -527 -792 -522
rect -754 -527 -749 -522
rect -810 -547 -805 -542
rect -672 -547 -667 -542
rect -795 -557 -790 -552
rect -446 -464 -441 -459
rect -411 -461 -406 -456
rect -752 -568 -747 -563
rect -639 -591 -635 -587
rect -639 -613 -635 -609
rect -367 -474 -362 -469
rect -411 -614 -407 -610
rect -190 -575 -185 -570
rect -127 -474 -122 -469
rect -91 -475 -86 -470
rect -71 -475 -66 -470
rect -34 -498 -29 -493
rect 45 -505 50 -500
rect -143 -526 -138 -521
rect -106 -526 -100 -520
rect -91 -527 -86 -522
rect -48 -527 -43 -522
rect 34 -547 39 -542
rect -89 -557 -84 -552
rect -46 -568 -41 -563
rect -190 -611 -185 -606
rect -734 -624 -729 -619
rect 42 -624 47 -619
rect -556 -639 -551 -634
rect 40 -639 45 -634
rect -377 -659 -372 -654
rect -7 -659 -2 -654
rect -165 -675 -160 -670
rect 94 -675 101 -670
rect -970 -737 -965 -732
rect -734 -713 -729 -708
rect -675 -713 -671 -709
rect -556 -713 -551 -708
rect -497 -713 -492 -708
rect -376 -713 -371 -708
rect -317 -713 -313 -709
rect -165 -713 -160 -708
rect -748 -721 -743 -716
rect -909 -737 -904 -732
rect -570 -721 -565 -716
rect -390 -721 -385 -716
rect -179 -721 -174 -716
rect -106 -714 -101 -707
rect -866 -792 -861 -787
rect -411 -800 -406 -795
rect -561 -807 -557 -803
rect -974 -923 -969 -918
rect -708 -876 -703 -871
rect -683 -876 -678 -871
rect -661 -876 -655 -870
rect -678 -887 -673 -882
rect -482 -876 -477 -871
rect -457 -876 -452 -871
rect -422 -875 -417 -870
rect -447 -887 -442 -882
rect -264 -876 -259 -871
rect -239 -876 -234 -871
rect -619 -911 -614 -906
rect -401 -911 -396 -906
rect -831 -924 -826 -919
rect -422 -944 -417 -939
rect -447 -950 -442 -945
rect -660 -1081 -655 -1076
rect -401 -947 -396 -942
rect -225 -978 -220 -973
rect -79 -866 -74 -861
rect -70 -874 -65 -869
rect 53 -889 58 -884
rect -106 -944 -101 -939
rect -72 -945 -67 -940
rect -52 -945 -47 -940
rect -15 -968 -10 -963
rect 62 -975 67 -970
rect -207 -996 -202 -991
rect -190 -996 -185 -991
rect -87 -996 -81 -990
rect -72 -997 -67 -992
rect -29 -997 -24 -992
rect 53 -1017 58 -1012
rect -70 -1027 -65 -1022
rect -27 -1038 -22 -1033
rect -207 -1070 -203 -1066
rect -660 -1114 -655 -1109
rect -422 -1114 -417 -1109
rect -207 -1114 -203 -1110
rect 84 -1089 88 -1085
rect -734 -1129 -729 -1124
rect 42 -1129 47 -1124
rect -556 -1144 -551 -1139
rect 40 -1144 45 -1139
rect -377 -1164 -372 -1159
rect -7 -1164 -2 -1159
rect 84 -1170 88 -1166
rect 141 -158 146 -153
rect 141 -659 146 -654
rect 187 -139 192 -134
rect 187 -639 192 -634
rect 303 -80 308 -75
rect 371 -80 376 -75
rect 247 -118 252 -113
rect 285 -505 290 -500
rect 248 -624 253 -619
rect 330 -568 335 -563
rect 331 -639 336 -634
rect 285 -681 290 -676
rect 331 -1068 336 -1063
rect 259 -1105 264 -1100
rect 299 -1105 304 -1100
rect 331 -1124 336 -1119
rect 248 -1129 253 -1124
rect 187 -1144 192 -1139
rect 141 -1164 146 -1159
rect -165 -1180 -160 -1175
rect 94 -1180 101 -1175
rect -974 -1242 -969 -1237
rect -734 -1218 -729 -1213
rect -675 -1218 -670 -1213
rect -556 -1218 -551 -1213
rect -497 -1218 -492 -1213
rect -376 -1218 -371 -1213
rect -317 -1218 -313 -1214
rect -165 -1218 -160 -1213
rect -106 -1218 -102 -1214
rect -748 -1226 -743 -1221
rect -920 -1242 -915 -1237
rect -570 -1226 -565 -1221
rect -390 -1226 -385 -1221
rect -179 -1226 -174 -1221
rect -660 -1318 -656 -1314
rect -831 -1350 -826 -1345
rect -422 -1337 -418 -1333
rect -753 -1441 -748 -1436
rect -728 -1441 -723 -1436
rect -693 -1440 -688 -1435
rect -724 -1452 -719 -1447
rect -527 -1441 -522 -1436
rect -502 -1441 -497 -1436
rect -469 -1440 -464 -1435
rect -492 -1452 -487 -1447
rect -309 -1441 -304 -1436
rect -284 -1441 -279 -1436
rect -242 -1440 -237 -1435
rect -892 -1476 -888 -1472
rect -664 -1476 -659 -1471
rect -446 -1476 -441 -1471
rect -725 -1513 -720 -1508
rect -693 -1513 -688 -1508
rect -645 -1510 -640 -1505
rect -423 -1510 -418 -1505
rect -79 -1430 -74 -1425
rect -70 -1438 -65 -1433
rect 53 -1453 58 -1448
rect -270 -1510 -265 -1505
rect -106 -1508 -101 -1503
rect -72 -1509 -67 -1504
rect -52 -1509 -47 -1504
rect -15 -1532 -10 -1527
rect 62 -1539 67 -1534
rect -207 -1561 -202 -1556
rect -87 -1560 -81 -1554
rect -72 -1561 -67 -1556
rect -29 -1561 -24 -1556
rect 53 -1581 58 -1576
rect -70 -1591 -65 -1586
rect -27 -1602 -22 -1597
rect -446 -1617 -442 -1613
<< pm12contact >>
rect -564 -420 -559 -415
rect -501 -420 -496 -415
rect -532 -429 -527 -424
rect -477 -428 -472 -423
rect -312 -420 -307 -415
rect -249 -420 -244 -415
rect -280 -429 -275 -424
rect -225 -428 -220 -423
rect -786 -890 -781 -885
rect -723 -890 -718 -885
rect -754 -899 -749 -894
rect -699 -898 -694 -893
rect -560 -890 -555 -885
rect -497 -890 -492 -885
rect -528 -899 -523 -894
rect -473 -898 -468 -893
rect -342 -890 -337 -885
rect -279 -890 -274 -885
rect -310 -899 -305 -894
rect -255 -898 -250 -893
rect -831 -1455 -826 -1450
rect -768 -1455 -763 -1450
rect -799 -1464 -794 -1459
rect -744 -1463 -739 -1458
rect -605 -1455 -600 -1450
rect -542 -1455 -537 -1450
rect -573 -1464 -568 -1459
rect -518 -1463 -513 -1458
rect -387 -1455 -382 -1450
rect -324 -1455 -319 -1450
rect -355 -1464 -350 -1459
rect -300 -1463 -295 -1458
<< metal2 >>
rect -28 127 -24 128
rect -364 123 403 127
rect -364 -12 -360 123
rect -350 -4 -345 101
rect -990 -33 -923 -29
rect -283 -56 -279 -9
rect -242 -12 -238 123
rect -228 -4 -223 79
rect -159 -41 -155 -9
rect -128 -12 -124 123
rect -114 -4 -109 58
rect -49 -41 -45 -9
rect -28 -12 -24 123
rect -14 -4 -9 36
rect 69 -9 335 -5
rect -558 -60 -279 -56
rect -960 -251 -931 -247
rect -846 -275 -576 -271
rect -972 -547 -898 -543
rect -965 -737 -909 -733
rect -866 -787 -862 -336
rect -846 -485 -842 -275
rect -558 -295 -554 -60
rect -463 -80 303 -76
rect -463 -230 -459 -80
rect -449 -222 -444 -118
rect -379 -271 -375 -227
rect -533 -275 -375 -271
rect -332 -283 -328 -92
rect -305 -230 -301 -80
rect -291 -222 -286 -139
rect -232 -293 -228 -227
rect -166 -230 -162 -80
rect -152 -222 -147 -158
rect -564 -298 -554 -295
rect -540 -297 -228 -293
rect -564 -302 -560 -298
rect -646 -390 -642 -336
rect -803 -458 -800 -396
rect -812 -461 -800 -458
rect -812 -520 -809 -461
rect -795 -470 -792 -404
rect -795 -473 -777 -470
rect -795 -484 -792 -473
rect -795 -493 -792 -489
rect -795 -496 -740 -493
rect -846 -547 -810 -543
rect -795 -552 -792 -527
rect -752 -563 -749 -527
rect -670 -542 -667 -419
rect -540 -416 -536 -297
rect -92 -313 -88 -227
rect -288 -317 -88 -313
rect -481 -405 -461 -401
rect -559 -420 -501 -416
rect -527 -428 -477 -424
rect -623 -479 -619 -441
rect -446 -459 -442 -417
rect -411 -456 -407 -405
rect -288 -416 -284 -317
rect -74 -326 -70 -95
rect -48 -230 -44 -80
rect 68 -118 247 -113
rect 70 -139 187 -134
rect 63 -158 141 -153
rect -34 -181 95 -176
rect -34 -222 -29 -181
rect -143 -330 -70 -326
rect -229 -405 -209 -401
rect -307 -420 -249 -416
rect -275 -428 -225 -424
rect -367 -469 -363 -442
rect -204 -479 -200 -417
rect -623 -483 -200 -479
rect -658 -505 -635 -501
rect -639 -587 -635 -505
rect -190 -570 -186 -405
rect -143 -521 -139 -330
rect 56 -347 60 -227
rect -127 -351 60 -347
rect -127 -469 -123 -351
rect -97 -458 -94 -396
rect -106 -461 -94 -458
rect -106 -520 -103 -461
rect -89 -470 -86 -404
rect -86 -473 -71 -470
rect -89 -493 -86 -475
rect -89 -496 -34 -493
rect -89 -552 -86 -527
rect -46 -563 -43 -527
rect 36 -542 39 -419
rect 50 -505 285 -501
rect 331 -563 335 -9
rect 376 -80 400 -76
rect -748 -600 413 -596
rect -748 -716 -744 -600
rect -570 -601 -557 -600
rect -734 -708 -729 -624
rect -675 -809 -671 -713
rect -639 -803 -635 -613
rect -570 -716 -566 -601
rect -556 -708 -551 -639
rect -639 -807 -561 -803
rect -762 -813 -671 -809
rect -762 -886 -758 -813
rect -497 -818 -493 -713
rect -411 -795 -407 -614
rect -390 -716 -386 -600
rect -376 -708 -371 -659
rect -317 -816 -313 -713
rect -536 -822 -493 -818
rect -318 -820 -313 -816
rect -703 -875 -683 -871
rect -781 -890 -723 -886
rect -749 -898 -699 -894
rect -969 -923 -831 -919
rect -678 -1066 -674 -887
rect -831 -1070 -674 -1066
rect -969 -1242 -920 -1238
rect -831 -1345 -827 -1070
rect -660 -1076 -656 -876
rect -536 -886 -532 -822
rect -477 -875 -457 -871
rect -555 -890 -497 -886
rect -523 -898 -473 -894
rect -619 -968 -615 -911
rect -447 -945 -443 -887
rect -422 -939 -418 -875
rect -318 -886 -314 -820
rect -259 -875 -239 -871
rect -337 -890 -279 -886
rect -305 -898 -255 -894
rect -401 -942 -397 -911
rect -619 -972 -269 -968
rect -273 -1062 -269 -972
rect -225 -1062 -221 -978
rect -190 -991 -186 -611
rect -179 -716 -175 -600
rect 47 -624 248 -619
rect 45 -639 187 -634
rect -2 -659 141 -654
rect -165 -708 -160 -675
rect -106 -939 -102 -714
rect -78 -928 -75 -866
rect -87 -931 -75 -928
rect -87 -990 -84 -931
rect -70 -940 -67 -874
rect -67 -943 -52 -940
rect -70 -963 -67 -945
rect -70 -966 -15 -963
rect -273 -1066 -221 -1062
rect -207 -1066 -203 -996
rect -70 -1022 -67 -997
rect -27 -1033 -24 -997
rect 55 -1012 58 -889
rect 67 -975 88 -971
rect 84 -1085 88 -975
rect -748 -1105 259 -1101
rect -748 -1221 -744 -1105
rect -570 -1106 -557 -1105
rect -734 -1213 -729 -1129
rect -675 -1358 -671 -1218
rect -660 -1314 -656 -1114
rect -570 -1221 -566 -1106
rect -556 -1213 -551 -1144
rect -497 -1346 -493 -1218
rect -422 -1333 -418 -1114
rect -390 -1221 -386 -1105
rect -376 -1213 -371 -1164
rect -317 -1259 -313 -1218
rect -363 -1263 -313 -1259
rect -807 -1362 -671 -1358
rect -581 -1350 -493 -1346
rect -807 -1451 -803 -1362
rect -748 -1440 -728 -1436
rect -826 -1455 -768 -1451
rect -794 -1463 -744 -1459
rect -892 -1535 -888 -1476
rect -724 -1508 -720 -1452
rect -693 -1508 -689 -1440
rect -581 -1451 -577 -1350
rect -522 -1440 -502 -1436
rect -600 -1455 -542 -1451
rect -568 -1463 -518 -1459
rect -664 -1506 -660 -1476
rect -664 -1510 -645 -1506
rect -492 -1535 -488 -1452
rect -892 -1539 -488 -1535
rect -469 -1694 -465 -1440
rect -363 -1451 -359 -1263
rect -304 -1440 -284 -1436
rect -382 -1455 -324 -1451
rect -350 -1463 -300 -1459
rect -446 -1613 -442 -1476
rect -418 -1510 -270 -1506
rect -242 -1699 -238 -1440
rect -207 -1556 -203 -1114
rect -179 -1221 -175 -1105
rect 47 -1129 248 -1124
rect 45 -1144 187 -1139
rect -2 -1164 141 -1159
rect -165 -1213 -160 -1180
rect -106 -1503 -102 -1218
rect 84 -1379 88 -1170
rect 84 -1383 142 -1379
rect -78 -1492 -75 -1430
rect -87 -1495 -75 -1492
rect -87 -1554 -84 -1495
rect -70 -1504 -67 -1438
rect -67 -1507 -52 -1504
rect -70 -1527 -67 -1509
rect -70 -1530 -15 -1527
rect -70 -1586 -67 -1561
rect -27 -1597 -24 -1561
rect 55 -1576 58 -1453
rect 67 -1539 97 -1535
rect 93 -1699 97 -1539
rect 138 -1699 142 -1383
rect 285 -1699 289 -681
rect 331 -1063 335 -639
rect 331 -1070 335 -1068
rect 304 -1105 382 -1101
rect 331 -1699 335 -1124
<< labels >>
rlabel metal1 -951 17 -946 21 1 VDD
rlabel metal1 -918 -33 -910 -29 1 GND
rlabel metal2 396 123 403 127 5 A0
rlabel metal1 267 101 273 106 1 B3
rlabel metal1 211 79 217 84 1 B2
rlabel metal1 153 58 159 63 1 B1
rlabel metal1 112 36 118 41 1 B0
rlabel metal2 393 -80 400 -76 1 A1
rlabel metal2 406 -600 413 -596 7 A2
rlabel metal2 376 -1105 382 -1101 1 A3
rlabel metal2 331 -1699 335 -1694 1 S0
rlabel metal2 285 -1699 289 -1694 1 S1
rlabel metal2 138 -1699 142 -1694 1 S2
rlabel metal2 93 -1699 97 -1694 1 S3
rlabel metal2 -242 -1699 -238 -1694 1 S4
rlabel metal2 -469 -1694 -465 -1689 1 S5
rlabel metal1 -693 -1699 -689 -1694 1 S6
rlabel metal1 -724 -1699 -720 -1694 1 C
<< end >>
