magic
tech scmos
timestamp 1667580020
<< nwell >>
rect -24 -5 26 19
<< ntransistor >>
rect 13 -18 15 -14
rect -13 -27 -11 -23
rect -3 -27 -1 -23
<< ptransistor >>
rect -13 1 -11 9
rect -3 1 -1 9
rect 13 1 15 9
<< ndiffusion >>
rect 12 -18 13 -14
rect 15 -18 16 -14
rect -14 -27 -13 -23
rect -11 -27 -3 -23
rect -1 -27 0 -23
<< pdiffusion >>
rect -14 1 -13 9
rect -11 1 -8 9
rect -4 1 -3 9
rect -1 1 0 9
rect 12 1 13 9
rect 15 1 16 9
<< ndcontact >>
rect 8 -18 12 -14
rect 16 -18 20 -14
rect -18 -27 -14 -23
rect 0 -27 4 -23
<< pdcontact >>
rect -18 1 -14 9
rect -8 1 -4 9
rect 0 1 4 9
rect 8 1 12 9
rect 16 1 20 9
<< polysilicon >>
rect -13 9 -11 12
rect -3 9 -1 12
rect 13 9 15 12
rect -13 -23 -11 1
rect -3 -23 -1 1
rect 13 -14 15 1
rect -13 -30 -11 -27
rect -3 -30 -1 -27
rect 13 -30 15 -18
<< polycontact >>
rect -17 -11 -13 -7
rect -7 -19 -3 -15
rect 9 -11 13 -7
<< metal1 >>
rect -24 15 26 19
rect -18 9 -14 15
rect 0 9 4 15
rect 8 9 12 15
rect -8 -2 -4 1
rect -8 -5 4 -2
rect 0 -7 4 -5
rect 16 -7 20 1
rect -19 -11 -17 -7
rect 0 -11 9 -7
rect 16 -11 26 -7
rect -19 -19 -7 -15
rect 0 -23 4 -11
rect 16 -14 20 -11
rect -18 -31 -14 -27
rect 8 -31 12 -18
rect -24 -35 26 -31
<< labels >>
rlabel metal1 -18 -9 -18 -9 1 A
rlabel metal1 -1 18 -1 18 5 VDD
rlabel metal1 -18 -17 -18 -17 1 B
rlabel metal1 -1 -34 -1 -34 1 GND
rlabel metal1 23 -9 23 -9 7 C
rlabel metal1 6 -9 6 -9 1 node1
<< end >>
