magic
tech scmos
timestamp 1667649636
<< nwell >>
rect 6 -223 56 -203
rect -51 -303 -27 -283
rect -9 -303 47 -283
rect -51 -355 -27 -335
<< ntransistor >>
rect 43 -236 45 -232
rect 17 -245 19 -241
rect 27 -245 29 -241
rect -40 -315 -38 -311
rect -40 -367 -38 -363
rect 4 -367 6 -363
rect 13 -367 15 -363
rect 22 -367 24 -363
rect 32 -367 34 -363
<< ptransistor >>
rect 17 -217 19 -209
rect 27 -217 29 -209
rect 43 -217 45 -209
rect -40 -297 -38 -289
rect 3 -297 5 -289
rect 13 -297 15 -289
rect 23 -297 25 -289
rect 32 -297 34 -289
rect -40 -349 -38 -341
<< ndiffusion >>
rect 42 -236 43 -232
rect 45 -236 46 -232
rect 16 -245 17 -241
rect 19 -245 27 -241
rect 29 -245 30 -241
rect -41 -315 -40 -311
rect -38 -315 -37 -311
rect -41 -367 -40 -363
rect -38 -367 -37 -363
rect 2 -367 4 -363
rect 6 -367 13 -363
rect 15 -367 17 -363
rect 21 -367 22 -363
rect 24 -367 32 -363
rect 34 -367 35 -363
<< pdiffusion >>
rect 16 -217 17 -209
rect 19 -217 22 -209
rect 26 -217 27 -209
rect 29 -217 30 -209
rect 42 -217 43 -209
rect 45 -217 46 -209
rect -41 -297 -40 -289
rect -38 -297 -37 -289
rect 1 -297 3 -289
rect 5 -297 13 -289
rect 15 -297 17 -289
rect 21 -297 23 -289
rect 25 -297 32 -289
rect 34 -297 35 -289
rect -41 -349 -40 -341
rect -38 -349 -37 -341
<< ndcontact >>
rect 38 -236 42 -232
rect 46 -236 50 -232
rect 12 -245 16 -241
rect 30 -245 34 -241
rect -45 -315 -41 -311
rect -37 -315 -33 -311
rect -45 -367 -41 -363
rect -37 -367 -33 -363
rect -3 -367 2 -363
rect 17 -367 21 -363
rect 35 -367 39 -363
<< pdcontact >>
rect 12 -217 16 -209
rect 22 -217 26 -209
rect 30 -217 34 -209
rect 38 -217 42 -209
rect 46 -217 50 -209
rect -45 -297 -41 -289
rect -37 -297 -33 -289
rect -3 -297 1 -289
rect 17 -297 21 -289
rect 35 -297 39 -289
rect -45 -349 -41 -341
rect -37 -349 -33 -341
<< polysilicon >>
rect 17 -209 19 -206
rect 27 -209 29 -206
rect 43 -209 45 -206
rect 17 -241 19 -217
rect 27 -241 29 -217
rect 43 -232 45 -217
rect 17 -248 19 -245
rect 27 -248 29 -245
rect 43 -248 45 -236
rect 3 -279 43 -277
rect -40 -289 -38 -286
rect 3 -289 5 -279
rect 13 -289 15 -286
rect 23 -289 25 -286
rect 32 -289 34 -286
rect -40 -311 -38 -297
rect 3 -308 5 -297
rect -40 -318 -38 -315
rect 13 -319 15 -297
rect -3 -321 15 -319
rect -40 -341 -38 -338
rect -3 -344 -1 -321
rect 23 -326 25 -297
rect 13 -328 25 -326
rect -3 -346 6 -344
rect -40 -363 -38 -349
rect 4 -363 6 -346
rect 13 -363 15 -328
rect 32 -346 34 -297
rect 22 -348 34 -346
rect 22 -363 24 -348
rect 41 -353 43 -279
rect 32 -355 43 -353
rect 32 -363 34 -355
rect -40 -370 -38 -367
rect 4 -391 6 -367
rect 13 -371 15 -367
rect 22 -402 24 -367
rect 32 -371 34 -367
<< polycontact >>
rect 13 -229 17 -225
rect 23 -237 27 -233
rect 39 -229 43 -225
rect -44 -308 -40 -304
rect -1 -308 3 -304
rect 9 -331 13 -327
rect -44 -360 -40 -356
rect 0 -391 4 -387
rect 18 -402 22 -398
<< metal1 >>
rect -87 -203 56 -200
rect -87 -279 -83 -203
rect 12 -209 16 -203
rect 30 -209 34 -203
rect 38 -209 42 -203
rect 22 -220 26 -217
rect 22 -223 34 -220
rect 30 -225 34 -223
rect 46 -225 50 -217
rect -75 -229 13 -225
rect 30 -229 39 -225
rect 46 -229 56 -225
rect -66 -237 23 -233
rect 30 -241 34 -229
rect 46 -232 50 -229
rect 12 -249 16 -245
rect 38 -249 42 -236
rect 6 -253 52 -249
rect -87 -283 49 -279
rect -95 -308 -73 -304
rect -60 -331 -56 -283
rect -45 -289 -41 -283
rect -3 -289 1 -283
rect 35 -289 39 -283
rect -37 -304 -33 -297
rect -48 -308 -44 -304
rect -37 -308 -1 -304
rect -37 -311 -33 -308
rect -45 -321 -41 -315
rect -48 -325 -20 -321
rect -60 -335 -27 -331
rect -45 -341 -41 -335
rect -24 -344 -20 -325
rect -11 -331 9 -327
rect 17 -335 21 -297
rect 17 -339 52 -335
rect -24 -348 -10 -344
rect -95 -360 -88 -356
rect -37 -356 -33 -349
rect -82 -360 -73 -356
rect -68 -360 -44 -356
rect -37 -360 -30 -356
rect -37 -363 -33 -360
rect -45 -377 -41 -367
rect -14 -377 -10 -348
rect 17 -363 21 -339
rect -3 -377 2 -367
rect 35 -377 39 -367
rect -86 -381 52 -377
rect -66 -391 0 -387
rect -23 -402 18 -398
<< m2contact >>
rect -80 -230 -75 -225
rect -71 -238 -66 -233
rect 52 -253 57 -248
rect -73 -309 -68 -304
rect -53 -309 -48 -304
rect -16 -332 -11 -327
rect -88 -360 -82 -354
rect -73 -361 -68 -356
rect -30 -361 -25 -356
rect 52 -381 57 -376
rect -71 -391 -66 -386
rect -28 -402 -23 -397
<< metal2 >>
rect -79 -292 -76 -230
rect -88 -295 -76 -292
rect -88 -354 -85 -295
rect -71 -304 -68 -238
rect -68 -307 -53 -304
rect -71 -327 -68 -309
rect -71 -330 -16 -327
rect -71 -386 -68 -361
rect -28 -397 -25 -361
rect 54 -376 57 -253
<< labels >>
rlabel metal1 48 -339 52 -335 7 SUM
rlabel metal1 -86 -381 49 -377 1 GND
rlabel metal1 -86 -283 49 -279 1 VDD
rlabel metal1 36 -227 36 -227 1 node1
rlabel metal1 -95 -308 -91 -304 3 A
rlabel metal1 -95 -360 -91 -356 3 B
rlabel metal1 52 -229 56 -225 7 CARRY
<< end >>
