*** FULL ADDER

.INCLUDE ../TSMC_180nm.txt
.INCLUDE ../MULTIPLIER/INVERTER.sub

*PARAMETERS
.PARAM X=90nm

.PARAM Width_p=4*X
.PARAM Length_p=2*X

.PARAM Width_n=2*X
.PARAM Length_n=2*X

.PARAM supply=1
.global gnd vdd

.temp 25

*NET-LIST

*FULL ADDER

*CARRY
*  -------------------------------------------------------VDD
*          |           |                   | 
*   A -- |Mp1|   B --|Mp2|          B -- |Mp4|    
*          |           |                   | 
*          -------------                   |-------node3
*                |                         |
*                ---------node1     A -- |Mp5|
*                |                         |
*         ---- |Mp3|                       |         _____
*    C____|      |_________________________|_________CARRY____|inverter|___CARRY     
*         |      |                         |
*         ---- |Mn3|                       |
*                |                         |
*                ---------node2     A -- |Mn5|
*                |                         |
*          -------------                   |-------node4
*          |           |                   |    
*   A -- |Mn1|   B --|Mn2|          B -- |Mn4|     
*          |           |                   | 
* -------------------------------------------------------GND   

*SUM
*--------------------------------------------------------VDD
*         |            |            |              |
*  A -- |Mp6|   B -- |Mp7|   C -- |Mp8|     A -- |Mp10|
*         |____________|____________|              |______node7
*                      |                           |
*                      ---------node5       B -- |Mp11|
*                      |                           |______node8
*               -----|Mp9|                         |
*              |       |                    C -- |Mp12|
*     _____    |       |                           |              ___
*     CARRY ---        -------------------------------------------SUM---|inverter|----SUM
*              |       |                           |
*              |       |                    C -- |Mn12|
*               -----|Mn9|                         |______node9
*                      |                           |
*                      ---------node6        B -- |Mn11|
*         _____________|____________               |______node10 
*         |            |            |              |
*  A -- |Mn6|   B -- |Mn7|   C -- |Mn8|     A -- |Mn10|
*         |            |            |              |
*--------------------------------------------------------GND
*
Mp1 node1  A  vdd  vdd CMOSP W={2*Width_p} L={Length_p}
Mp2 node1  B  vdd  vdd CMOSP W={2*Width_p} L={Length_p}
Mp3 CARRY_ C node1 vdd CMOSP W={2*Width_p} L={Length_p}

Mn1 node2  A  gnd  gnd CMOSN W={2*Width_n} L={Length_n}
Mn2 node2  B  gnd  gnd CMOSN W={2*Width_n} L={Length_n}
Mn3 CARRY_ C node2 gnd CMOSN W={2*Width_n} L={Length_n}

Mp4 node3  B  vdd  vdd CMOSP W={2*Width_p} L={Length_p}
Mp5 CARRY_ A node3 vdd CMOSP W={2*Width_p} L={Length_p}

Mn4 node4  B  gnd  gnd CMOSN W={2*Width_n} L={Length_n}
Mn5 CARRY_ A node4 gnd CMOSN W={2*Width_n} L={Length_n}

xinv1 CARRY_ vdd gnd CARRY INVERTER

Mp6 node5  A      vdd   vdd CMOSP W={2*Width_p} L={Length_p}
Mp7 node5  B      vdd   vdd CMOSP W={2*Width_p} L={Length_p}
Mp8 node5  C      vdd   vdd CMOSP W={2*Width_p} L={Length_p}
Mp9 SUM_  CARRY_ node5  vdd CMOSP W={2*Width_p} L={Length_p}

Mn6 node6  A      gnd   gnd CMOSN W={2*Width_n} L={Length_n}
Mn7 node6  A      gnd   gnd CMOSN W={2*Width_n} L={Length_n}
Mn8 node6  A      gnd   gnd CMOSN W={2*Width_n} L={Length_n}
Mn9 SUM_  CARRY_ node6  gnd CMOSN W={2*Width_n} L={Length_n}

Mp10 node7  A   vdd   vdd CMOSP W={2*Width_p} L={Length_p}
Mp11 node8  B  node7  vdd CMOSP W={2*Width_p} L={Length_p}
Mp12 SUM_   C  node8  vdd CMOSP W={2*Width_p} L={Length_p}

Mn10 node10 A   gnd   gnd CMOSN W={2*Width_n} L={Length_n}
Mn11 node 9 B  node10 gnd CMOSN W={2*Width_n} L={Length_n}
Mn12 SUM_   C  node9  gnd CMOSN W={2*Width_n} L={Length_n}

xinv2 SUM_ vdd gnd SUM INVERTER

*SOURCE
VDD vdd gnd 'supply'

*Capacitive LOAD
CL1 SUM gnd 2f
CL2 CARRY gnd 2f

*INPUT WAVEFORM
VinA A gnd 0
VinB B gnd 0
VinC c gnd 0

*ANALYSIS
.op

*CONTROL COMMANDS
.CONTROL
    alter VinA = 0
    alter VinB = 0
    alter VinC = 0
    op
    let leakage_power = -1*VDD#branch+(v(A)*(-VinA#branch))+(v(B)*(-VinB#branch))+(v(C)*(-VinC#branch))
    echo "VA = 0 VB = 0 VC = 0">>"FA_Pre_Layout_leakage.txt"
    echo "Leakage Power = $&leakage_power">>"FA_Pre_Layout_leakage.txt"

    alter VinA = 0
    alter VinB = 0
    alter VinC = 1
    op
    let leakage_power = -1*VDD#branch+(v(A)*(-VinA#branch))+(v(B)*(-VinB#branch))+(v(C)*(-VinC#branch))
    echo "VA = 0 VB = 0 VC = 1">>"FA_Pre_Layout_leakage.txt"
    echo "Leakage Power = $&leakage_power">>"FA_Pre_Layout_leakage.txt"

    alter VinA = 0
    alter VinB = 1
    alter VinC = 0
    op
    let leakage_power = -1*VDD#branch+(v(A)*(-VinA#branch))+(v(B)*(-VinB#branch))+(v(C)*(-VinC#branch))
    echo "VA = 0 VB = 1 VC = 0">>"FA_Pre_Layout_leakage.txt"
    echo "Leakage Power = $&leakage_power">>"FA_Pre_Layout_leakage.txt"

    alter VinA = 0
    alter VinB = 1
    alter VinC = 1
    op
    let leakage_power = -1*VDD#branch+(v(A)*(-VinA#branch))+(v(B)*(-VinB#branch))+(v(C)*(-VinC#branch))
    echo "VA = 0 VB = 1 VC = 1">>"FA_Pre_Layout_leakage.txt"
    echo "Leakage Power = $&leakage_power">>"FA_Pre_Layout_leakage.txt"

    alter VinA = 1
    alter VinB = 0
    alter VinC = 0
    op
    let leakage_power = -1*VDD#branch+(v(A)*(-VinA#branch))+(v(B)*(-VinB#branch))+(v(C)*(-VinC#branch))
    echo "VA = 1 VB = 0 VC = 0">>"FA_Pre_Layout_leakage.txt"
    echo "Leakage Power = $&leakage_power">>"FA_Pre_Layout_leakage.txt"

    alter VinA = 1
    alter VinB = 0
    alter VinC = 1
    op
    let leakage_power = -1*VDD#branch+(v(A)*(-VinA#branch))+(v(B)*(-VinB#branch))+(v(C)*(-VinC#branch))
    echo "VA = 1 VB = 0 VC = 1">>"FA_Pre_Layout_leakage.txt"
    echo "Leakage Power = $&leakage_power">>"FA_Pre_Layout_leakage.txt"

    alter VinA = 1
    alter VinB = 1
    alter VinC = 0
    op
    let leakage_power = -1*VDD#branch+(v(A)*(-VinA#branch))+(v(B)*(-VinB#branch))+(v(C)*(-VinC#branch))
    echo "VA = 1 VB = 1 VC = 0">>"FA_Pre_Layout_leakage.txt"
    echo "Leakage Power = $&leakage_power">>"FA_Pre_Layout_leakage.txt"

    alter VinA = 1
    alter VinB = 1
    alter VinC = 1
    op
    let leakage_power = -1*VDD#branch+(v(A)*(-VinA#branch))+(v(B)*(-VinB#branch))+(v(C)*(-VinC#branch))
    echo "VA = 1 VB = 1 VC = 1">>"FA_Pre_Layout_leakage.txt"
    echo "Leakage Power = $&leakage_power">>"FA_Pre_Layout_leakage.txt"


.ENDC
.END